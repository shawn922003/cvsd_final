module power_to_tuple_63_51(
    input  [5:0] i_power,
    output reg [5:0] o_tuple
);

    always @(*) begin
        case (i_power)
            6'd63: o_tuple = 6'b000000;  // ZERO (not in ALPHA_POLY_BITS)

            6'd0:  o_tuple = 6'b000001;  // alpha^0  = [1,0,0,0,0,0]  -> 000001
            6'd1:  o_tuple = 6'b000010;  // alpha^1
            6'd2:  o_tuple = 6'b000100;  // alpha^2
            6'd3:  o_tuple = 6'b001000;  // alpha^3
            6'd4:  o_tuple = 6'b010000;  // alpha^4
            6'd5:  o_tuple = 6'b100000;  // alpha^5
            6'd6:  o_tuple = 6'b000011;  // alpha^6
            6'd7:  o_tuple = 6'b000110;  // alpha^7
            6'd8:  o_tuple = 6'b001100;  // alpha^8
            6'd9:  o_tuple = 6'b011000;  // alpha^9
            6'd10: o_tuple = 6'b110000;  // alpha^10
            6'd11: o_tuple = 6'b100011;  // alpha^11
            6'd12: o_tuple = 6'b000101;  // alpha^12
            6'd13: o_tuple = 6'b001010;  // alpha^13
            6'd14: o_tuple = 6'b010100;  // alpha^14
            6'd15: o_tuple = 6'b101000;  // alpha^15
            6'd16: o_tuple = 6'b010011;  // alpha^16
            6'd17: o_tuple = 6'b100110;  // alpha^17
            6'd18: o_tuple = 6'b001111;  // alpha^18
            6'd19: o_tuple = 6'b011110;  // alpha^19
            6'd20: o_tuple = 6'b111100;  // alpha^20
            6'd21: o_tuple = 6'b111011;  // alpha^21
            6'd22: o_tuple = 6'b110101;  // alpha^22
            6'd23: o_tuple = 6'b101001;  // alpha^23
            6'd24: o_tuple = 6'b010001;  // alpha^24
            6'd25: o_tuple = 6'b100010;  // alpha^25
            6'd26: o_tuple = 6'b001110;  // alpha^26
            6'd27: o_tuple = 6'b011100;  // alpha^27
            6'd28: o_tuple = 6'b111000;  // alpha^28
            6'd29: o_tuple = 6'b110001;  // alpha^29
            6'd30: o_tuple = 6'b110011;  // alpha^30
            6'd31: o_tuple = 6'b100101;  // alpha^31
            6'd32: o_tuple = 6'b001001;  // alpha^32
            6'd33: o_tuple = 6'b010010;  // alpha^33
            6'd34: o_tuple = 6'b100100;  // alpha^34
            6'd35: o_tuple = 6'b001011;  // alpha^35
            6'd36: o_tuple = 6'b010110;  // alpha^36
            6'd37: o_tuple = 6'b101100;  // alpha^37
            6'd38: o_tuple = 6'b011011;  // alpha^38
            6'd39: o_tuple = 6'b110110;  // alpha^39
            6'd40: o_tuple = 6'b101111;  // alpha^40
            6'd41: o_tuple = 6'b011101;  // alpha^41
            6'd42: o_tuple = 6'b111010;  // alpha^42
            6'd43: o_tuple = 6'b110111;  // alpha^43
            6'd44: o_tuple = 6'b101011;  // alpha^44
            6'd45: o_tuple = 6'b011001;  // alpha^45
            6'd46: o_tuple = 6'b110010;  // alpha^46
            6'd47: o_tuple = 6'b100111;  // alpha^47
            6'd48: o_tuple = 6'b001101;  // alpha^48
            6'd49: o_tuple = 6'b011010;  // alpha^49
            6'd50: o_tuple = 6'b110100;  // alpha^50
            6'd51: o_tuple = 6'b101011;  // alpha^51
            6'd52: o_tuple = 6'b010101;  // alpha^52
            6'd53: o_tuple = 6'b101010;  // alpha^53
            6'd54: o_tuple = 6'b010111;  // alpha^54
            6'd55: o_tuple = 6'b101110;  // alpha^55
            6'd56: o_tuple = 6'b011111;  // alpha^56
            6'd57: o_tuple = 6'b111110;  // alpha^57
            6'd58: o_tuple = 6'b111111;  // alpha^58
            6'd59: o_tuple = 6'b111101;  // alpha^59
            6'd60: o_tuple = 6'b111001;  // alpha^60
            6'd61: o_tuple = 6'b110001;  // alpha^61
            6'd62: o_tuple = 6'b100001;  // alpha^62
        endcase
    end

endmodule


module tuple_to_power_63_51(
    input  [5:0] i_tuple,
    output reg [5:0] o_power
);

    always @(*) begin
        case (i_tuple)
            6'b000000: o_power = 6'd63;  // ZERO ( -1)

            6'b000001: o_power = 6'd0;   // alpha^0
            6'b000010: o_power = 6'd1;   // alpha^1
            6'b000100: o_power = 6'd2;   // alpha^2
            6'b001000: o_power = 6'd3;   // alpha^3
            6'b010000: o_power = 6'd4;   // alpha^4
            6'b100000: o_power = 6'd5;   // alpha^5
            6'b000011: o_power = 6'd6;   // alpha^6
            6'b000110: o_power = 6'd7;   // alpha^7
            6'b001100: o_power = 6'd8;   // alpha^8
            6'b011000: o_power = 6'd9;   // alpha^9
            6'b110000: o_power = 6'd10;  // alpha^10
            6'b100011: o_power = 6'd11;  // alpha^11
            6'b000101: o_power = 6'd12;  // alpha^12
            6'b001010: o_power = 6'd13;  // alpha^13
            6'b010100: o_power = 6'd14;  // alpha^14
            6'b101000: o_power = 6'd15;  // alpha^15
            6'b010011: o_power = 6'd16;  // alpha^16
            6'b100110: o_power = 6'd17;  // alpha^17
            6'b001111: o_power = 6'd18;  // alpha^18
            6'b011110: o_power = 6'd19;  // alpha^19
            6'b111100: o_power = 6'd20;  // alpha^20
            6'b111011: o_power = 6'd21;  // alpha^21
            6'b110101: o_power = 6'd22;  // alpha^22
            6'b101001: o_power = 6'd23;  // alpha^23
            6'b010001: o_power = 6'd24;  // alpha^24
            6'b100010: o_power = 6'd25;  // alpha^25
            6'b001110: o_power = 6'd26;  // alpha^26
            6'b011100: o_power = 6'd27;  // alpha^27
            6'b111000: o_power = 6'd28;  // alpha^28
            6'b110001: o_power = 6'd29;  // alpha^29
            6'b110011: o_power = 6'd30;  // alpha^30
            6'b100101: o_power = 6'd31;  // alpha^31
            6'b001001: o_power = 6'd32;  // alpha^32
            6'b010010: o_power = 6'd33;  // alpha^33
            6'b100100: o_power = 6'd34;  // alpha^34
            6'b001011: o_power = 6'd35;  // alpha^35
            6'b010110: o_power = 6'd36;  // alpha^36
            6'b101100: o_power = 6'd37;  // alpha^37
            6'b011011: o_power = 6'd38;  // alpha^38
            6'b110110: o_power = 6'd39;  // alpha^39
            6'b101111: o_power = 6'd40;  // alpha^40
            6'b011101: o_power = 6'd41;  // alpha^41
            6'b111010: o_power = 6'd42;  // alpha^42
            6'b110111: o_power = 6'd43;  // alpha^43
            6'b101011: o_power = 6'd44;  // alpha^44
            6'b011001: o_power = 6'd45;  // alpha^45
            6'b110010: o_power = 6'd46;  // alpha^46
            6'b100111: o_power = 6'd47;  // alpha^47
            6'b001101: o_power = 6'd48;  // alpha^48
            6'b011010: o_power = 6'd49;  // alpha^49
            6'b110100: o_power = 6'd50;  // alpha^50
            6'b101011: o_power = 6'd51;  // alpha^51
            6'b010101: o_power = 6'd52;  // alpha^52
            6'b101010: o_power = 6'd53;  // alpha^53
            6'b010111: o_power = 6'd54;  // alpha^54
            6'b101110: o_power = 6'd55;  // alpha^55
            6'b011111: o_power = 6'd56;  // alpha^56
            6'b111110: o_power = 6'd57;  // alpha^57
            6'b111111: o_power = 6'd58;  // alpha^58
            6'b111101: o_power = 6'd59;  // alpha^59
            6'b111001: o_power = 6'd60;  // alpha^60
            6'b110001: o_power = 6'd61;  // alpha^61
            6'b100001: o_power = 6'd62;  // alpha^62

        endcase
    end

endmodule





// BCH (255, 239) Galois Field GF(2^8) Lookup Tables
// Primitive polynomial: p(x) = 1 + x^2 + x^3 + x^4 + x^8
// Generated from Python bch_table.py

module power_to_tuple_255(
    input  [7:0] i_power,
    output reg [7:0] o_tuple
);

    always @(*) begin
        case (i_power)
            8'd255: o_tuple = 8'b00000000;  // ZERO
            8'd0:   o_tuple = 8'b00000001;  // [1,0,0,0,0,0,0,0]
            8'd1:   o_tuple = 8'b00000010;  // [0,1,0,0,0,0,0,0]
            8'd2:   o_tuple = 8'b00000100;  // [0,0,1,0,0,0,0,0]
            8'd3:   o_tuple = 8'b00001000;  // [0,0,0,1,0,0,0,0]
            8'd4:   o_tuple = 8'b00010000;  // [0,0,0,0,1,0,0,0]
            8'd5:   o_tuple = 8'b00100000;  // [0,0,0,0,0,1,0,0]
            8'd6:   o_tuple = 8'b01000000;  // [0,0,0,0,0,0,1,0]
            8'd7:   o_tuple = 8'b10000000;  // [0,0,0,0,0,0,0,1]
            8'd8:   o_tuple = 8'b00011101;  // [1,0,1,1,1,0,0,0]
            8'd9:   o_tuple = 8'b00111010;  // [0,1,0,1,1,1,0,0]
            8'd10:  o_tuple = 8'b01110100;  // [0,0,1,0,1,1,1,0]
            8'd11:  o_tuple = 8'b11101000;  // [0,0,0,1,0,1,1,1]
            8'd12:  o_tuple = 8'b11001101;  // [1,0,1,1,0,0,1,1]
            8'd13:  o_tuple = 8'b10010111;  // [1,1,1,0,1,0,0,1]
            8'd14:  o_tuple = 8'b00110011;  // [1,1,0,0,1,1,0,0]
            8'd15:  o_tuple = 8'b01100110;  // [0,1,1,0,0,1,1,0]
            8'd16:  o_tuple = 8'b11001100;  // [0,0,1,1,0,0,1,1]
            8'd17:  o_tuple = 8'b10000101;  // [1,0,1,0,0,0,0,1]
            8'd18:  o_tuple = 8'b00010111;  // [1,1,1,0,1,0,0,0]
            8'd19:  o_tuple = 8'b00101110;  // [0,1,1,1,0,1,0,0]
            8'd20:  o_tuple = 8'b01011100;  // [0,0,1,1,1,0,1,0]
            8'd21:  o_tuple = 8'b10111000;  // [0,0,0,1,1,1,0,1]
            8'd22:  o_tuple = 8'b01101101;  // [1,0,1,1,0,1,1,0]
            8'd23:  o_tuple = 8'b11011010;  // [0,1,0,1,1,0,1,1]
            8'd24:  o_tuple = 8'b10101001;  // [1,0,0,1,0,1,0,1]
            8'd25:  o_tuple = 8'b01001111;  // [1,1,1,1,0,0,1,0]
            8'd26:  o_tuple = 8'b10011110;  // [0,1,1,1,1,0,0,1]
            8'd27:  o_tuple = 8'b00110001;  // [1,0,0,0,1,1,0,0]
            8'd28:  o_tuple = 8'b01100010;  // [0,1,0,0,0,1,1,0]
            8'd29:  o_tuple = 8'b11000100;  // [0,0,1,0,0,0,1,1]
            8'd30:  o_tuple = 8'b10010101;  // [1,0,1,0,1,0,0,1]
            8'd31:  o_tuple = 8'b00110111;  // [1,1,1,0,1,1,0,0]
            8'd32:  o_tuple = 8'b01101110;  // [0,1,1,1,0,1,1,0]
            8'd33:  o_tuple = 8'b11011100;  // [0,0,1,1,1,0,1,1]
            8'd34:  o_tuple = 8'b10100101;  // [1,0,1,0,0,1,0,1]
            8'd35:  o_tuple = 8'b01010111;  // [1,1,1,0,1,0,1,0]
            8'd36:  o_tuple = 8'b10101110;  // [0,1,1,1,0,1,0,1]
            8'd37:  o_tuple = 8'b01000001;  // [1,0,0,0,0,0,1,0]
            8'd38:  o_tuple = 8'b10000010;  // [0,1,0,0,0,0,0,1]
            8'd39:  o_tuple = 8'b00011001;  // [1,0,0,1,1,0,0,0]
            8'd40:  o_tuple = 8'b00110010;  // [0,1,0,0,1,1,0,0]
            8'd41:  o_tuple = 8'b01100100;  // [0,0,1,0,0,1,1,0]
            8'd42:  o_tuple = 8'b11001000;  // [0,0,0,1,0,0,1,1]
            8'd43:  o_tuple = 8'b10001101;  // [1,0,1,1,0,0,0,1]
            8'd44:  o_tuple = 8'b00000111;  // [1,1,1,0,0,0,0,0]
            8'd45:  o_tuple = 8'b00001110;  // [0,1,1,1,0,0,0,0]
            8'd46:  o_tuple = 8'b00011100;  // [0,0,1,1,1,0,0,0]
            8'd47:  o_tuple = 8'b00111000;  // [0,0,0,1,1,1,0,0]
            8'd48:  o_tuple = 8'b01110000;  // [0,0,0,0,1,1,1,0]
            8'd49:  o_tuple = 8'b11100000;  // [0,0,0,0,0,1,1,1]
            8'd50:  o_tuple = 8'b11011101;  // [1,0,1,1,1,0,1,1]
            8'd51:  o_tuple = 8'b10100111;  // [1,1,1,0,0,1,0,1]
            8'd52:  o_tuple = 8'b01010011;  // [1,1,0,0,1,0,1,0]
            8'd53:  o_tuple = 8'b10100110;  // [0,1,1,0,0,1,0,1]
            8'd54:  o_tuple = 8'b01010001;  // [1,0,0,0,1,0,1,0]
            8'd55:  o_tuple = 8'b10100010;  // [0,1,0,0,0,1,0,1]
            8'd56:  o_tuple = 8'b01011001;  // [1,0,0,1,1,0,1,0]
            8'd57:  o_tuple = 8'b10110010;  // [0,1,0,0,1,1,0,1]
            8'd58:  o_tuple = 8'b01111001;  // [1,0,0,1,1,1,1,0]
            8'd59:  o_tuple = 8'b11110010;  // [0,1,0,0,1,1,1,1]
            8'd60:  o_tuple = 8'b11111001;  // [1,0,0,1,1,1,1,1]
            8'd61:  o_tuple = 8'b11101111;  // [1,1,1,1,0,1,1,1]
            8'd62:  o_tuple = 8'b11000011;  // [1,1,0,0,0,0,1,1]
            8'd63:  o_tuple = 8'b10011011;  // [1,1,0,1,1,0,0,1]
            8'd64:  o_tuple = 8'b00101011;  // [1,1,0,1,0,1,0,0]
            8'd65:  o_tuple = 8'b01010110;  // [0,1,1,0,1,0,1,0]
            8'd66:  o_tuple = 8'b10101100;  // [0,0,1,1,0,1,0,1]
            8'd67:  o_tuple = 8'b01000101;  // [1,0,1,0,0,0,1,0]
            8'd68:  o_tuple = 8'b10001010;  // [0,1,0,1,0,0,0,1]
            8'd69:  o_tuple = 8'b00001001;  // [1,0,0,1,0,0,0,0]
            8'd70:  o_tuple = 8'b00010010;  // [0,1,0,0,1,0,0,0]
            8'd71:  o_tuple = 8'b00100100;  // [0,0,1,0,0,1,0,0]
            8'd72:  o_tuple = 8'b01001000;  // [0,0,0,1,0,0,1,0]
            8'd73:  o_tuple = 8'b10010000;  // [0,0,0,0,1,0,0,1]
            8'd74:  o_tuple = 8'b00111101;  // [1,0,1,1,1,1,0,0]
            8'd75:  o_tuple = 8'b01111010;  // [0,1,0,1,1,1,1,0]
            8'd76:  o_tuple = 8'b11110100;  // [0,0,1,0,1,1,1,1]
            8'd77:  o_tuple = 8'b11110101;  // [1,0,1,0,1,1,1,1]
            8'd78:  o_tuple = 8'b11110111;  // [1,1,1,0,1,1,1,1]
            8'd79:  o_tuple = 8'b11110011;  // [1,1,0,0,1,1,1,1]
            8'd80:  o_tuple = 8'b11111011;  // [1,1,0,1,1,1,1,1]
            8'd81:  o_tuple = 8'b11101011;  // [1,1,0,1,0,1,1,1]
            8'd82:  o_tuple = 8'b11001011;  // [1,1,0,1,0,0,1,1]
            8'd83:  o_tuple = 8'b10001011;  // [1,1,0,1,0,0,0,1]
            8'd84:  o_tuple = 8'b00001011;  // [1,1,0,1,0,0,0,0]
            8'd85:  o_tuple = 8'b00010110;  // [0,1,1,0,1,0,0,0]
            8'd86:  o_tuple = 8'b00101100;  // [0,0,1,1,0,1,0,0]
            8'd87:  o_tuple = 8'b01011000;  // [0,0,0,1,1,0,1,0]
            8'd88:  o_tuple = 8'b10110000;  // [0,0,0,0,1,1,0,1]
            8'd89:  o_tuple = 8'b01111101;  // [1,0,1,1,1,1,1,0]
            8'd90:  o_tuple = 8'b11111010;  // [0,1,0,1,1,1,1,1]
            8'd91:  o_tuple = 8'b11101001;  // [1,0,0,1,0,1,1,1]
            8'd92:  o_tuple = 8'b11001111;  // [1,1,1,1,0,0,1,1]
            8'd93:  o_tuple = 8'b10010011;  // [1,1,0,0,1,0,0,1]
            8'd94:  o_tuple = 8'b00111011;  // [1,1,0,1,1,1,0,0]
            8'd95:  o_tuple = 8'b01110110;  // [0,1,1,0,1,1,1,0]
            8'd96:  o_tuple = 8'b11101100;  // [0,0,1,1,0,1,1,1]
            8'd97:  o_tuple = 8'b11000101;  // [1,0,1,0,0,0,1,1]
            8'd98:  o_tuple = 8'b10010111;  // [1,1,1,0,1,0,0,1]
            8'd99:  o_tuple = 8'b00110011;  // [1,1,0,0,1,1,0,0]
            8'd100: o_tuple = 8'b01100110;  // [0,1,1,0,0,1,1,0]
            8'd101: o_tuple = 8'b11001100;  // [0,0,1,1,0,0,1,1]
            8'd102: o_tuple = 8'b10000101;  // [1,0,1,0,0,0,0,1]
            8'd103: o_tuple = 8'b00010111;  // [1,1,1,0,1,0,0,0]
            8'd104: o_tuple = 8'b00101110;  // [0,1,1,1,0,1,0,0]
            8'd105: o_tuple = 8'b01011100;  // [0,0,1,1,1,0,1,0]
            8'd106: o_tuple = 8'b10111000;  // [0,0,0,1,1,1,0,1]
            8'd107: o_tuple = 8'b01101101;  // [1,0,1,1,0,1,1,0]
            8'd108: o_tuple = 8'b11011010;  // [0,1,0,1,1,0,1,1]
            8'd109: o_tuple = 8'b10101001;  // [1,0,0,1,0,1,0,1]
            8'd110: o_tuple = 8'b01001111;  // [1,1,1,1,0,0,1,0]
            8'd111: o_tuple = 8'b10011110;  // [0,1,1,1,1,0,0,1]
            8'd112: o_tuple = 8'b00110001;  // [1,0,0,0,1,1,0,0]
            8'd113: o_tuple = 8'b01100010;  // [0,1,0,0,0,1,1,0]
            8'd114: o_tuple = 8'b11000100;  // [0,0,1,0,0,0,1,1]
            8'd115: o_tuple = 8'b10010101;  // [1,0,1,0,1,0,0,1]
            8'd116: o_tuple = 8'b00110111;  // [1,1,1,0,1,1,0,0]
            8'd117: o_tuple = 8'b01101110;  // [0,1,1,1,0,1,1,0]
            8'd118: o_tuple = 8'b11011100;  // [0,0,1,1,1,0,1,1]
            8'd119: o_tuple = 8'b10100101;  // [1,0,1,0,0,1,0,1]
            8'd120: o_tuple = 8'b01010111;  // [1,1,1,0,1,0,1,0]
            8'd121: o_tuple = 8'b10101110;  // [0,1,1,1,0,1,0,1]
            8'd122: o_tuple = 8'b01000001;  // [1,0,0,0,0,0,1,0]
            8'd123: o_tuple = 8'b10000010;  // [0,1,0,0,0,0,0,1]
            8'd124: o_tuple = 8'b00011001;  // [1,0,0,1,1,0,0,0]
            8'd125: o_tuple = 8'b00110010;  // [0,1,0,0,1,1,0,0]
            8'd126: o_tuple = 8'b01100100;  // [0,0,1,0,0,1,1,0]
            8'd127: o_tuple = 8'b11001000;  // [0,0,0,1,0,0,1,1]
            8'd128: o_tuple = 8'b10001101;  // [1,0,1,1,0,0,0,1]
            8'd129: o_tuple = 8'b00000111;  // [1,1,1,0,0,0,0,0]
            8'd130: o_tuple = 8'b00001110;  // [0,1,1,1,0,0,0,0]
            8'd131: o_tuple = 8'b00011100;  // [0,0,1,1,1,0,0,0]
            8'd132: o_tuple = 8'b00111000;  // [0,0,0,1,1,1,0,0]
            8'd133: o_tuple = 8'b01110000;  // [0,0,0,0,1,1,1,0]
            8'd134: o_tuple = 8'b11100000;  // [0,0,0,0,0,1,1,1]
            8'd135: o_tuple = 8'b11011101;  // [1,0,1,1,1,0,1,1]
            8'd136: o_tuple = 8'b10100111;  // [1,1,1,0,0,1,0,1]
            8'd137: o_tuple = 8'b01010011;  // [1,1,0,0,1,0,1,0]
            8'd138: o_tuple = 8'b10100110;  // [0,1,1,0,0,1,0,1]
            8'd139: o_tuple = 8'b01010001;  // [1,0,0,0,1,0,1,0]
            8'd140: o_tuple = 8'b10100010;  // [0,1,0,0,0,1,0,1]
            8'd141: o_tuple = 8'b01011001;  // [1,0,0,1,1,0,1,0]
            8'd142: o_tuple = 8'b10110010;  // [0,1,0,0,1,1,0,1]
            8'd143: o_tuple = 8'b01111001;  // [1,0,0,1,1,1,1,0]
            8'd144: o_tuple = 8'b11110010;  // [0,1,0,0,1,1,1,1]
            8'd145: o_tuple = 8'b11111001;  // [1,0,0,1,1,1,1,1]
            8'd146: o_tuple = 8'b11101111;  // [1,1,1,1,0,1,1,1]
            8'd147: o_tuple = 8'b11000011;  // [1,1,0,0,0,0,1,1]
            8'd148: o_tuple = 8'b10011011;  // [1,1,0,1,1,0,0,1]
            8'd149: o_tuple = 8'b00101011;  // [1,1,0,1,0,1,0,0]
            8'd150: o_tuple = 8'b01010110;  // [0,1,1,0,1,0,1,0]
            8'd151: o_tuple = 8'b10101100;  // [0,0,1,1,0,1,0,1]
            8'd152: o_tuple = 8'b01000101;  // [1,0,1,0,0,0,1,0]
            8'd153: o_tuple = 8'b10001010;  // [0,1,0,1,0,0,0,1]
            8'd154: o_tuple = 8'b00001001;  // [1,0,0,1,0,0,0,0]
            8'd155: o_tuple = 8'b00010010;  // [0,1,0,0,1,0,0,0]
            8'd156: o_tuple = 8'b00100100;  // [0,0,1,0,0,1,0,0]
            8'd157: o_tuple = 8'b01001000;  // [0,0,0,1,0,0,1,0]
            8'd158: o_tuple = 8'b10010000;  // [0,0,0,0,1,0,0,1]
            8'd159: o_tuple = 8'b00111101;  // [1,0,1,1,1,1,0,0]
            8'd160: o_tuple = 8'b01111010;  // [0,1,0,1,1,1,1,0]
            8'd161: o_tuple = 8'b11110100;  // [0,0,1,0,1,1,1,1]
            8'd162: o_tuple = 8'b11110101;  // [1,0,1,0,1,1,1,1]
            8'd163: o_tuple = 8'b11110111;  // [1,1,1,0,1,1,1,1]
            8'd164: o_tuple = 8'b11110011;  // [1,1,0,0,1,1,1,1]
            8'd165: o_tuple = 8'b11111011;  // [1,1,0,1,1,1,1,1]
            8'd166: o_tuple = 8'b11101011;  // [1,1,0,1,0,1,1,1]
            8'd167: o_tuple = 8'b11001011;  // [1,1,0,1,0,0,1,1]
            8'd168: o_tuple = 8'b10001011;  // [1,1,0,1,0,0,0,1]
            8'd169: o_tuple = 8'b00001011;  // [1,1,0,1,0,0,0,0]
            8'd170: o_tuple = 8'b00010110;  // [0,1,1,0,1,0,0,0]
            8'd171: o_tuple = 8'b00101100;  // [0,0,1,1,0,1,0,0]
            8'd172: o_tuple = 8'b01011000;  // [0,0,0,1,1,0,1,0]
            8'd173: o_tuple = 8'b10110000;  // [0,0,0,0,1,1,0,1]
            8'd174: o_tuple = 8'b01111101;  // [1,0,1,1,1,1,1,0]
            8'd175: o_tuple = 8'b11111010;  // [0,1,0,1,1,1,1,1]
            8'd176: o_tuple = 8'b11101001;  // [1,0,0,1,0,1,1,1]
            8'd177: o_tuple = 8'b11001111;  // [1,1,1,1,0,0,1,1]
            8'd178: o_tuple = 8'b10010011;  // [1,1,0,0,1,0,0,1]
            8'd179: o_tuple = 8'b00111011;  // [1,1,0,1,1,1,0,0]
            8'd180: o_tuple = 8'b01110110;  // [0,1,1,0,1,1,1,0]
            8'd181: o_tuple = 8'b11101100;  // [0,0,1,1,0,1,1,1]
            8'd182: o_tuple = 8'b11000101;  // [1,0,1,0,0,0,1,1]
            8'd183: o_tuple = 8'b10010111;  // [1,1,1,0,1,0,0,1]
            8'd184: o_tuple = 8'b00110011;  // [1,1,0,0,1,1,0,0]
            8'd185: o_tuple = 8'b01100110;  // [0,1,1,0,0,1,1,0]
            8'd186: o_tuple = 8'b11001100;  // [0,0,1,1,0,0,1,1]
            8'd187: o_tuple = 8'b10000101;  // [1,0,1,0,0,0,0,1]
            8'd188: o_tuple = 8'b00010111;  // [1,1,1,0,1,0,0,0]
            8'd189: o_tuple = 8'b00101110;  // [0,1,1,1,0,1,0,0]
            8'd190: o_tuple = 8'b01011100;  // [0,0,1,1,1,0,1,0]
            8'd191: o_tuple = 8'b10111000;  // [0,0,0,1,1,1,0,1]
            8'd192: o_tuple = 8'b01101101;  // [1,0,1,1,0,1,1,0]
            8'd193: o_tuple = 8'b11011010;  // [0,1,0,1,1,0,1,1]
            8'd194: o_tuple = 8'b10101001;  // [1,0,0,1,0,1,0,1]
            8'd195: o_tuple = 8'b01001111;  // [1,1,1,1,0,0,1,0]
            8'd196: o_tuple = 8'b10011110;  // [0,1,1,1,1,0,0,1]
            8'd197: o_tuple = 8'b00110001;  // [1,0,0,0,1,1,0,0]
            8'd198: o_tuple = 8'b01100010;  // [0,1,0,0,0,1,1,0]
            8'd199: o_tuple = 8'b11000100;  // [0,0,1,0,0,0,1,1]
            8'd200: o_tuple = 8'b10010101;  // [1,0,1,0,1,0,0,1]
            8'd201: o_tuple = 8'b00110111;  // [1,1,1,0,1,1,0,0]
            8'd202: o_tuple = 8'b01101110;  // [0,1,1,1,0,1,1,0]
            8'd203: o_tuple = 8'b11011100;  // [0,0,1,1,1,0,1,1]
            8'd204: o_tuple = 8'b10100101;  // [1,0,1,0,0,1,0,1]
            8'd205: o_tuple = 8'b01010111;  // [1,1,1,0,1,0,1,0]
            8'd206: o_tuple = 8'b10101110;  // [0,1,1,1,0,1,0,1]
            8'd207: o_tuple = 8'b01000001;  // [1,0,0,0,0,0,1,0]
            8'd208: o_tuple = 8'b10000010;  // [0,1,0,0,0,0,0,1]
            8'd209: o_tuple = 8'b00011001;  // [1,0,0,1,1,0,0,0]
            8'd210: o_tuple = 8'b00110010;  // [0,1,0,0,1,1,0,0]
            8'd211: o_tuple = 8'b01100100;  // [0,0,1,0,0,1,1,0]
            8'd212: o_tuple = 8'b11001000;  // [0,0,0,1,0,0,1,1]
            8'd213: o_tuple = 8'b10001101;  // [1,0,1,1,0,0,0,1]
            8'd214: o_tuple = 8'b00000111;  // [1,1,1,0,0,0,0,0]
            8'd215: o_tuple = 8'b00001110;  // [0,1,1,1,0,0,0,0]
            8'd216: o_tuple = 8'b00011100;  // [0,0,1,1,1,0,0,0]
            8'd217: o_tuple = 8'b00111000;  // [0,0,0,1,1,1,0,0]
            8'd218: o_tuple = 8'b01110000;  // [0,0,0,0,1,1,1,0]
            8'd219: o_tuple = 8'b11100000;  // [0,0,0,0,0,1,1,1]
            8'd220: o_tuple = 8'b11011101;  // [1,0,1,1,1,0,1,1]
            8'd221: o_tuple = 8'b10100111;  // [1,1,1,0,0,1,0,1]
            8'd222: o_tuple = 8'b01010011;  // [1,1,0,0,1,0,1,0]
            8'd223: o_tuple = 8'b10100110;  // [0,1,1,0,0,1,0,1]
            8'd224: o_tuple = 8'b01010001;  // [1,0,0,0,1,0,1,0]
            8'd225: o_tuple = 8'b10100010;  // [0,1,0,0,0,1,0,1]
            8'd226: o_tuple = 8'b01011001;  // [1,0,0,1,1,0,1,0]
            8'd227: o_tuple = 8'b10110010;  // [0,1,0,0,1,1,0,1]
            8'd228: o_tuple = 8'b01111001;  // [1,0,0,1,1,1,1,0]
            8'd229: o_tuple = 8'b11110010;  // [0,1,0,0,1,1,1,1]
            8'd230: o_tuple = 8'b11111001;  // [1,0,0,1,1,1,1,1]
            8'd231: o_tuple = 8'b11101111;  // [1,1,1,1,0,1,1,1]
            8'd232: o_tuple = 8'b11000011;  // [1,1,0,0,0,0,1,1]
            8'd233: o_tuple = 8'b10011011;  // [1,1,0,1,1,0,0,1]
            8'd234: o_tuple = 8'b00101011;  // [1,1,0,1,0,1,0,0]
            8'd235: o_tuple = 8'b01010110;  // [0,1,1,0,1,0,1,0]
            8'd236: o_tuple = 8'b10101100;  // [0,0,1,1,0,1,0,1]
            8'd237: o_tuple = 8'b01000101;  // [1,0,1,0,0,0,1,0]
            8'd238: o_tuple = 8'b10001010;  // [0,1,0,1,0,0,0,1]
            8'd239: o_tuple = 8'b00001001;  // [1,0,0,1,0,0,0,0]
            8'd240: o_tuple = 8'b00010010;  // [0,1,0,0,1,0,0,0]
            8'd241: o_tuple = 8'b00100100;  // [0,0,1,0,0,1,0,0]
            8'd242: o_tuple = 8'b01001000;  // [0,0,0,1,0,0,1,0]
            8'd243: o_tuple = 8'b10010000;  // [0,0,0,0,1,0,0,1]
            8'd244: o_tuple = 8'b00111101;  // [1,0,1,1,1,1,0,0]
            8'd245: o_tuple = 8'b01111010;  // [0,1,0,1,1,1,1,0]
            8'd246: o_tuple = 8'b11110100;  // [0,0,1,0,1,1,1,1]
            8'd247: o_tuple = 8'b11110101;  // [1,0,1,0,1,1,1,1]
            8'd248: o_tuple = 8'b11110111;  // [1,1,1,0,1,1,1,1]
            8'd249: o_tuple = 8'b11110011;  // [1,1,0,0,1,1,1,1]
            8'd250: o_tuple = 8'b11111011;  // [1,1,0,1,1,1,1,1]
            8'd251: o_tuple = 8'b11101011;  // [1,1,0,1,0,1,1,1]
            8'd252: o_tuple = 8'b11001011;  // [1,1,0,1,0,0,1,1]
            8'd253: o_tuple = 8'b10001011;  // [1,1,0,1,0,0,0,1]
            8'd254: o_tuple = 8'b00001011;  // [1,1,0,1,0,0,0,0]
            
            default: o_tuple = 8'b00000000;
        endcase
    end

endmodule


module tuple_to_power_255(
    input  [7:0] i_tuple,
    output reg [7:0] o_power
);

    always @(*) begin
        case (i_tuple)
            8'b00000000: o_power = 8'd255;  // ZERO
            8'b00000001: o_power = 8'd0;    // alpha^0
            8'b00000010: o_power = 8'd1;    // alpha^1
            8'b00000100: o_power = 8'd2;    // alpha^2
            8'b00001000: o_power = 8'd3;    // alpha^3
            8'b00010000: o_power = 8'd4;    // alpha^4
            8'b00100000: o_power = 8'd5;    // alpha^5
            8'b01000000: o_power = 8'd6;    // alpha^6
            8'b10000000: o_power = 8'd7;    // alpha^7
            8'b00011101: o_power = 8'd8;    // alpha^8
            8'b00111010: o_power = 8'd9;    // alpha^9
            8'b01110100: o_power = 8'd10;   // alpha^10
            8'b11101000: o_power = 8'd11;   // alpha^11
            8'b11001101: o_power = 8'd12;   // alpha^12
            8'b10110111: o_power = 8'd13;   // alpha^13
            8'b01110011: o_power = 8'd14;   // alpha^14
            8'b11100110: o_power = 8'd15;   // alpha^15
            8'b11110001: o_power = 8'd16;   // alpha^16
            8'b11111111: o_power = 8'd17;   // alpha^17
            8'b11101011: o_power = 8'd18;   // alpha^18
            8'b11001011: o_power = 8'd19;   // alpha^19
            8'b10101011: o_power = 8'd20;   // alpha^20
            8'b01101011: o_power = 8'd21;   // alpha^21
            8'b11010110: o_power = 8'd22;   // alpha^22
            8'b10010001: o_power = 8'd23;   // alpha^23
            8'b10101001: o_power = 8'd24;   // alpha^24
            8'b01001111: o_power = 8'd25;   // alpha^25
            8'b10011110: o_power = 8'd26;   // alpha^26
            8'b00110001: o_power = 8'd27;   // alpha^27
            8'b01100010: o_power = 8'd28;   // alpha^28
            8'b11000100: o_power = 8'd29;   // alpha^29
            8'b10010101: o_power = 8'd30;   // alpha^30
            8'b00110111: o_power = 8'd31;   // alpha^31
            8'b01101110: o_power = 8'd32;   // alpha^32
            8'b11011100: o_power = 8'd33;   // alpha^33
            8'b10100101: o_power = 8'd34;   // alpha^34
            8'b01010111: o_power = 8'd35;   // alpha^35
            8'b10101110: o_power = 8'd36;   // alpha^36
            8'b01000001: o_power = 8'd37;   // alpha^37
            8'b10000010: o_power = 8'd38;   // alpha^38
            8'b00011001: o_power = 8'd39;   // alpha^39
            8'b00110010: o_power = 8'd40;   // alpha^40
            8'b01100100: o_power = 8'd41;   // alpha^41
            8'b11001000: o_power = 8'd42;   // alpha^42
            8'b10001101: o_power = 8'd43;   // alpha^43
            8'b00000111: o_power = 8'd44;   // alpha^44
            8'b00001110: o_power = 8'd45;   // alpha^45
            8'b00011100: o_power = 8'd46;   // alpha^46
            8'b00111000: o_power = 8'd47;   // alpha^47
            8'b01110000: o_power = 8'd48;   // alpha^48
            8'b11100000: o_power = 8'd49;   // alpha^49
            8'b11011101: o_power = 8'd50;   // alpha^50
            8'b10100111: o_power = 8'd51;   // alpha^51
            8'b01010011: o_power = 8'd52;   // alpha^52
            8'b10100110: o_power = 8'd53;   // alpha^53
            8'b01010001: o_power = 8'd54;   // alpha^54
            8'b10100010: o_power = 8'd55;   // alpha^55
            8'b01011001: o_power = 8'd56;   // alpha^56
            8'b10110010: o_power = 8'd57;   // alpha^57
            8'b01111001: o_power = 8'd58;   // alpha^58
            8'b11110010: o_power = 8'd59;   // alpha^59
            8'b11111001: o_power = 8'd60;   // alpha^60
            8'b11101111: o_power = 8'd61;   // alpha^61
            8'b11000011: o_power = 8'd62;   // alpha^62
            8'b10011011: o_power = 8'd63;   // alpha^63
            8'b00101011: o_power = 8'd64;   // alpha^64
            8'b01010110: o_power = 8'd65;   // alpha^65
            8'b10101100: o_power = 8'd66;   // alpha^66
            8'b01000101: o_power = 8'd67;   // alpha^67
            8'b10001010: o_power = 8'd68;   // alpha^68
            8'b00001001: o_power = 8'd69;   // alpha^69
            8'b00010010: o_power = 8'd70;   // alpha^70
            8'b00100100: o_power = 8'd71;   // alpha^71
            8'b01001000: o_power = 8'd72;   // alpha^72
            8'b10010000: o_power = 8'd73;   // alpha^73
            8'b00111101: o_power = 8'd74;   // alpha^74
            8'b01111010: o_power = 8'd75;   // alpha^75
            8'b11110100: o_power = 8'd76;   // alpha^76
            8'b11110101: o_power = 8'd77;   // alpha^77
            8'b11110111: o_power = 8'd78;   // alpha^78
            8'b11110011: o_power = 8'd79;   // alpha^79
            8'b11111011: o_power = 8'd80;   // alpha^80
            8'b10001011: o_power = 8'd83;   // alpha^83
            8'b00001011: o_power = 8'd84;   // alpha^84
            8'b00010110: o_power = 8'd85;   // alpha^85
            8'b00101100: o_power = 8'd86;   // alpha^86
            8'b01011000: o_power = 8'd87;   // alpha^87
            8'b10110000: o_power = 8'd88;   // alpha^88
            8'b01111101: o_power = 8'd89;   // alpha^89
            8'b11111010: o_power = 8'd90;   // alpha^90
            8'b11101001: o_power = 8'd91;   // alpha^91
            8'b11001111: o_power = 8'd92;   // alpha^92
            8'b10010011: o_power = 8'd93;   // alpha^93
            8'b00111011: o_power = 8'd94;   // alpha^94
            8'b01110110: o_power = 8'd95;   // alpha^95
            8'b11101100: o_power = 8'd96;   // alpha^96
            8'b11000101: o_power = 8'd97;   // alpha^97
            8'b10010111: o_power = 8'd98;   // alpha^98
            8'b00110011: o_power = 8'd99;   // alpha^99
            8'b01100110: o_power = 8'd100;  // alpha^100
            8'b11001100: o_power = 8'd101;  // alpha^101
            8'b10000101: o_power = 8'd102;  // alpha^102
            8'b00010111: o_power = 8'd103;  // alpha^103
            8'b00101110: o_power = 8'd104;  // alpha^104
            8'b01011100: o_power = 8'd105;  // alpha^105
            8'b10111000: o_power = 8'd106;  // alpha^106
            8'b01101101: o_power = 8'd107;  // alpha^107
            8'b11011010: o_power = 8'd108;  // alpha^108
            8'b10101001: o_power = 8'd109;  // alpha^109
            8'b01001111: o_power = 8'd110;  // alpha^110
            8'b10011110: o_power = 8'd111;  // alpha^111
            8'b00110001: o_power = 8'd112;  // alpha^112
            8'b01100010: o_power = 8'd113;  // alpha^113
            8'b11000100: o_power = 8'd114;  // alpha^114
            8'b10010101: o_power = 8'd115;  // alpha^115
            8'b00110111: o_power = 8'd116;  // alpha^116
            8'b01101110: o_power = 8'd117;  // alpha^117
            8'b11011100: o_power = 8'd118;  // alpha^118
            8'b10100101: o_power = 8'd119;   // alpha^119
            8'b01010111: o_power = 8'd120;   // alpha^120
            8'b10101110: o_power = 8'd121;   // alpha^121
            8'b01000001: o_power = 8'd122;   // alpha^122
            8'b10000010: o_power = 8'd123;   // alpha^123
            8'b00011001: o_power = 8'd124;   // alpha^124
            8'b00110010: o_power = 8'd125;   // alpha^125
            8'b01100100: o_power = 8'd126;   // alpha^126
            8'b11001000: o_power = 8'd127;   // alpha^127
            8'b10001101: o_power = 8'd128;   // alpha^128
            8'b00000111: o_power = 8'd129;   // alpha^129
            8'b00001110: o_power = 8'd130;   // alpha^130
            8'b00011100: o_power = 8'd131;   // alpha^131
            8'b00111000: o_power = 8'd132;   // alpha^132
            8'b01110000: o_power = 8'd133;   // alpha^133
            8'b11100000: o_power = 8'd134;   // alpha^134
            8'b11011101: o_power = 8'd135;   // alpha^135
            8'b10100111: o_power = 8'd136;   // alpha^136
            8'b01010011: o_power = 8'd137;   // alpha^137
            8'b10100110: o_power = 8'd138;   // alpha^138
            8'b01010001: o_power = 8'd139;   // alpha^139
            8'b10100010: o_power = 8'd140;   // alpha^140
            8'b01011001: o_power = 8'd141;   // alpha^141
            8'b10110010: o_power = 8'd142;   // alpha^142
            8'b01111001: o_power = 8'd143;   // alpha^143
            8'b11110010: o_power = 8'd144;   // alpha^144
            8'b11111001: o_power = 8'd145;   // alpha^145
            8'b11101111: o_power = 8'd146;   // alpha^146
            8'b11000011: o_power = 8'd147;   // alpha^147
            8'b10011011: o_power = 8'd148;   // alpha^148
            8'b00101011: o_power = 8'd149;   // alpha^149
            8'b01010110: o_power = 8'd150;   // alpha^150
            8'b10101100: o_power = 8'd151;   // alpha^151
            8'b01000101: o_power = 8'd152;   // alpha^152
            8'b10001010: o_power = 8'd153;   // alpha^153
            8'b00001001: o_power = 8'd154;   // alpha^154
            8'b00010010: o_power = 8'd155;   // alpha^155
            8'b00100100: o_power = 8'd156;   // alpha^156
            8'b01001000: o_power = 8'd157;   // alpha^157
            8'b10010000: o_power = 8'd158;   // alpha^158
            8'b00111101: o_power = 8'd159;   // alpha^159
            8'b01111010: o_power = 8'd160;   // alpha^160
            8'b11110100: o_power = 8'd161;   // alpha^161
            8'b11110101: o_power = 8'd162;   // alpha^162
            8'b11110111: o_power = 8'd163;   // alpha^163
            8'b11110011: o_power = 8'd164;   // alpha^164
            8'b11111011: o_power = 8'd165;   // alpha^165
            8'b11101011: o_power = 8'd166;   // alpha^166
            8'b11001011: o_power = 8'd167;   // alpha^167
            8'b10001011: o_power = 8'd168;   // alpha^168
            8'b00001011: o_power = 8'd169;   // alpha^169
            8'b00010110: o_power = 8'd170;   // alpha^170
            8'b00101100: o_power = 8'd171;   // alpha^171
            8'b01011000: o_power = 8'd172;   // alpha^172
            8'b10110000: o_power = 8'd173;   // alpha^173
            8'b01111101: o_power = 8'd174;   // alpha^174
            8'b11111010: o_power = 8'd175;   // alpha^175
            8'b11101001: o_power = 8'd176;   // alpha^176
            8'b11001111: o_power = 8'd177;   // alpha^177
            8'b10010011: o_power = 8'd178;   // alpha^178
            8'b00111011: o_power = 8'd179;   // alpha^179
            8'b01110110: o_power = 8'd180;   // alpha^180
            8'b11101100: o_power = 8'd181;   // alpha^181
            8'b11000101: o_power = 8'd182;   // alpha^182
            8'b10010111: o_power = 8'd183;   // alpha^183
            8'b00110011: o_power = 8'd184;   // alpha^184
            8'b01100110: o_power = 8'd185;   // alpha^185
            8'b11001100: o_power = 8'd186;   // alpha^186
            8'b10000101: o_power = 8'd187;   // alpha^187
            8'b00010111: o_power = 8'd188;   // alpha^188
            8'b00101110: o_power = 8'd189;   // alpha^189
            8'b01011100: o_power = 8'd190;   // alpha^190
            8'b10111000: o_power = 8'd191;   // alpha^191
            8'b01101101: o_power = 8'd192;   // alpha^192
            8'b11011010: o_power = 8'd193;   // alpha^193
            8'b10101001: o_power = 8'd194;   // alpha^194
            8'b01001111: o_power = 8'd195;   // alpha^195
            8'b10011110: o_power = 8'd196;   // alpha^196
            8'b00110001: o_power = 8'd197;   // alpha^197
            8'b01100010: o_power = 8'd198;   // alpha^198
            8'b11000100: o_power = 8'd199;   // alpha^199
            8'b10010101: o_power = 8'd200;   // alpha^200
            8'b00110111: o_power = 8'd201;   // alpha^201
            8'b01101110: o_power = 8'd202;   // alpha^202
            8'b11011100: o_power = 8'd203;   // alpha^203
            8'b10100101: o_power = 8'd204;   // alpha^204
            8'b01010111: o_power = 8'd205;   // alpha^205
            8'b10101110: o_power = 8'd206;   // alpha^206
            8'b01000001: o_power = 8'd207;   // alpha^207
            8'b10000010: o_power = 8'd208;   // alpha^208
            8'b00011001: o_power = 8'd209;   // alpha^209
            8'b00110010: o_power = 8'd210;   // alpha^210
            8'b01100100: o_power = 8'd211;   // alpha^211
            8'b11001000: o_power = 8'd212;   // alpha^212
            8'b10001101: o_power = 8'd213;   // alpha^213
            8'b00000111: o_power = 8'd214;   // alpha^214
            8'b00001110: o_power = 8'd215;   // alpha^215
            8'b00011100: o_power = 8'd216;   // alpha^216
            8'b00111000: o_power = 8'd217;   // alpha^217
            8'b01110000: o_power = 8'd218;   // alpha^218
            8'b11100000: o_power = 8'd219;   // alpha^219
            8'b11011101: o_power = 8'd220;   // alpha^220
            8'b10100111: o_power = 8'd221;   // alpha^221
            8'b01010011: o_power = 8'd222;   // alpha^222
            8'b10100110: o_power = 8'd223;   // alpha^223
            8'b01010001: o_power = 8'd224;   // alpha^224
            8'b10100010: o_power = 8'd225;   // alpha^225
            8'b01011001: o_power = 8'd226;   // alpha^226
            8'b10110010: o_power = 8'd227;   // alpha^227
            8'b01111001: o_power = 8'd228;   // alpha^228
            8'b11110010: o_power = 8'd229;   // alpha^229
            8'b11111001: o_power = 8'd230;   // alpha^230
            8'b11101111: o_power = 8'd231;   // alpha^231
            8'b11000011: o_power = 8'd232;   // alpha^232
            8'b10011011: o_power = 8'd233;   // alpha^233
            8'b00101011: o_power = 8'd234;   // alpha^234
            8'b01010110: o_power = 8'd235;   // alpha^235
            8'b10101100: o_power = 8'd236;   // alpha^236
            8'b01000101: o_power = 8'd237;   // alpha^237
            8'b10001010: o_power = 8'd238;   // alpha^238
            8'b00001001: o_power = 8'd239;   // alpha^239
            8'b00010010: o_power = 8'd240;   // alpha^240
            8'b00100100: o_power = 8'd241;   // alpha^241
            8'b01001000: o_power = 8'd242;   // alpha^242
            8'b10010000: o_power = 8'd243;   // alpha^243
            8'b00111101: o_power = 8'd244;   // alpha^244
            8'b01111010: o_power = 8'd245;   // alpha^245
            8'b11110100: o_power = 8'd246;   // alpha^246
            8'b11110101: o_power = 8'd247;   // alpha^247
            8'b11110111: o_power = 8'd248;   // alpha^248
            8'b11110011: o_power = 8'd249;   // alpha^249
            8'b11111011: o_power = 8'd250;   // alpha^250
            8'b11101011: o_power = 8'd251;   // alpha^251
            8'b11001011: o_power = 8'd252;   // alpha^252
            8'b10001011: o_power = 8'd253;   // alpha^253
            8'b00001011: o_power = 8'd254;   // alpha^254 
            default: o_power = 8'd255;
        endcase
    end

endmodule




module power_to_tuple_1023_1015(
    input  [9:0] i_power,
    output reg [9:0] o_tuple
);

    always @(*) begin
        case (i_power)
            10'd1023: o_tuple = 10'b0000000000;  // ZERO (not in ALPHA_POLY_BITS)

            10'd   0: o_tuple = 10'b0000000001;  // alpha^0
            10'd   1: o_tuple = 10'b0000000010;  // alpha^1
            10'd   2: o_tuple = 10'b0000000100;  // alpha^2
            10'd   3: o_tuple = 10'b0000001000;  // alpha^3
            10'd   4: o_tuple = 10'b0000010000;  // alpha^4
            10'd   5: o_tuple = 10'b0000100000;  // alpha^5
            10'd   6: o_tuple = 10'b0001000000;  // alpha^6
            10'd   7: o_tuple = 10'b0010000000;  // alpha^7
            10'd   8: o_tuple = 10'b0100000000;  // alpha^8
            10'd   9: o_tuple = 10'b1000000000;  // alpha^9
            10'd  10: o_tuple = 10'b0000001001;  // alpha^10
            10'd  11: o_tuple = 10'b0000010010;  // alpha^11
            10'd  12: o_tuple = 10'b0000100100;  // alpha^12
            10'd  13: o_tuple = 10'b0001001000;  // alpha^13
            10'd  14: o_tuple = 10'b0010010000;  // alpha^14
            10'd  15: o_tuple = 10'b0100100000;  // alpha^15
            10'd  16: o_tuple = 10'b1001000000;  // alpha^16
            10'd  17: o_tuple = 10'b0010001001;  // alpha^17
            10'd  18: o_tuple = 10'b0100010010;  // alpha^18
            10'd  19: o_tuple = 10'b1000100100;  // alpha^19
            10'd  20: o_tuple = 10'b0001000001;  // alpha^20
            10'd  21: o_tuple = 10'b0010000010;  // alpha^21
            10'd  22: o_tuple = 10'b0100000100;  // alpha^22
            10'd  23: o_tuple = 10'b1000001000;  // alpha^23
            10'd  24: o_tuple = 10'b0000011001;  // alpha^24
            10'd  25: o_tuple = 10'b0000110010;  // alpha^25
            10'd  26: o_tuple = 10'b0001100100;  // alpha^26
            10'd  27: o_tuple = 10'b0011001000;  // alpha^27
            10'd  28: o_tuple = 10'b0110010000;  // alpha^28
            10'd  29: o_tuple = 10'b1100100000;  // alpha^29
            10'd  30: o_tuple = 10'b1001001001;  // alpha^30
            10'd  31: o_tuple = 10'b0010011011;  // alpha^31
            10'd  32: o_tuple = 10'b0100110110;  // alpha^32
            10'd  33: o_tuple = 10'b1001101100;  // alpha^33
            10'd  34: o_tuple = 10'b0011010001;  // alpha^34
            10'd  35: o_tuple = 10'b0110100010;  // alpha^35
            10'd  36: o_tuple = 10'b1101000100;  // alpha^36
            10'd  37: o_tuple = 10'b1010000001;  // alpha^37
            10'd  38: o_tuple = 10'b0100001011;  // alpha^38
            10'd  39: o_tuple = 10'b1000010110;  // alpha^39
            10'd  40: o_tuple = 10'b0000100101;  // alpha^40
            10'd  41: o_tuple = 10'b0001001010;  // alpha^41
            10'd  42: o_tuple = 10'b0010010100;  // alpha^42
            10'd  43: o_tuple = 10'b0100101000;  // alpha^43
            10'd  44: o_tuple = 10'b1001010000;  // alpha^44
            10'd  45: o_tuple = 10'b0010101001;  // alpha^45
            10'd  46: o_tuple = 10'b0101010010;  // alpha^46
            10'd  47: o_tuple = 10'b1010100100;  // alpha^47
            10'd  48: o_tuple = 10'b0101000001;  // alpha^48
            10'd  49: o_tuple = 10'b1010000010;  // alpha^49
            10'd  50: o_tuple = 10'b0100001101;  // alpha^50
            10'd  51: o_tuple = 10'b1000011010;  // alpha^51
            10'd  52: o_tuple = 10'b0000111101;  // alpha^52
            10'd  53: o_tuple = 10'b0001111010;  // alpha^53
            10'd  54: o_tuple = 10'b0011110100;  // alpha^54
            10'd  55: o_tuple = 10'b0111101000;  // alpha^55
            10'd  56: o_tuple = 10'b1111010000;  // alpha^56
            10'd  57: o_tuple = 10'b1110101001;  // alpha^57
            10'd  58: o_tuple = 10'b1101011011;  // alpha^58
            10'd  59: o_tuple = 10'b1010111111;  // alpha^59
            10'd  60: o_tuple = 10'b0101110111;  // alpha^60
            10'd  61: o_tuple = 10'b1011101110;  // alpha^61
            10'd  62: o_tuple = 10'b0111010101;  // alpha^62
            10'd  63: o_tuple = 10'b1110101010;  // alpha^63
            10'd  64: o_tuple = 10'b1101011101;  // alpha^64
            10'd  65: o_tuple = 10'b1010110011;  // alpha^65
            10'd  66: o_tuple = 10'b0101101111;  // alpha^66
            10'd  67: o_tuple = 10'b1011011110;  // alpha^67
            10'd  68: o_tuple = 10'b0110110101;  // alpha^68
            10'd  69: o_tuple = 10'b1101101010;  // alpha^69
            10'd  70: o_tuple = 10'b1011011101;  // alpha^70
            10'd  71: o_tuple = 10'b0110110011;  // alpha^71
            10'd  72: o_tuple = 10'b1101100110;  // alpha^72
            10'd  73: o_tuple = 10'b1011000101;  // alpha^73
            10'd  74: o_tuple = 10'b0110000011;  // alpha^74
            10'd  75: o_tuple = 10'b1100000110;  // alpha^75
            10'd  76: o_tuple = 10'b1000000101;  // alpha^76
            10'd  77: o_tuple = 10'b0000000011;  // alpha^77
            10'd  78: o_tuple = 10'b0000000110;  // alpha^78
            10'd  79: o_tuple = 10'b0000001100;  // alpha^79
            10'd  80: o_tuple = 10'b0000011000;  // alpha^80
            10'd  81: o_tuple = 10'b0000110000;  // alpha^81
            10'd  82: o_tuple = 10'b0001100000;  // alpha^82
            10'd  83: o_tuple = 10'b0011000000;  // alpha^83
            10'd  84: o_tuple = 10'b0110000000;  // alpha^84
            10'd  85: o_tuple = 10'b1100000000;  // alpha^85
            10'd  86: o_tuple = 10'b1000001001;  // alpha^86
            10'd  87: o_tuple = 10'b0000011011;  // alpha^87
            10'd  88: o_tuple = 10'b0000110110;  // alpha^88
            10'd  89: o_tuple = 10'b0001101100;  // alpha^89
            10'd  90: o_tuple = 10'b0011011000;  // alpha^90
            10'd  91: o_tuple = 10'b0110110000;  // alpha^91
            10'd  92: o_tuple = 10'b1101100000;  // alpha^92
            10'd  93: o_tuple = 10'b1011001001;  // alpha^93
            10'd  94: o_tuple = 10'b0110011011;  // alpha^94
            10'd  95: o_tuple = 10'b1100110110;  // alpha^95
            10'd  96: o_tuple = 10'b1001100101;  // alpha^96
            10'd  97: o_tuple = 10'b0011000011;  // alpha^97
            10'd  98: o_tuple = 10'b0110000110;  // alpha^98
            10'd  99: o_tuple = 10'b1100001100;  // alpha^99
            10'd 100: o_tuple = 10'b1000010001;  // alpha^100
            10'd 101: o_tuple = 10'b0000101011;  // alpha^101
            10'd 102: o_tuple = 10'b0001010110;  // alpha^102
            10'd 103: o_tuple = 10'b0010101100;  // alpha^103
            10'd 104: o_tuple = 10'b0101011000;  // alpha^104
            10'd 105: o_tuple = 10'b1010110000;  // alpha^105
            10'd 106: o_tuple = 10'b0101101001;  // alpha^106
            10'd 107: o_tuple = 10'b1011010010;  // alpha^107
            10'd 108: o_tuple = 10'b0110101101;  // alpha^108
            10'd 109: o_tuple = 10'b1101011010;  // alpha^109
            10'd 110: o_tuple = 10'b1010111101;  // alpha^110
            10'd 111: o_tuple = 10'b0101110011;  // alpha^111
            10'd 112: o_tuple = 10'b1011100110;  // alpha^112
            10'd 113: o_tuple = 10'b0111000101;  // alpha^113
            10'd 114: o_tuple = 10'b1110001010;  // alpha^114
            10'd 115: o_tuple = 10'b1100011101;  // alpha^115
            10'd 116: o_tuple = 10'b1000110011;  // alpha^116
            10'd 117: o_tuple = 10'b0001101111;  // alpha^117
            10'd 118: o_tuple = 10'b0011011110;  // alpha^118
            10'd 119: o_tuple = 10'b0110111100;  // alpha^119
            10'd 120: o_tuple = 10'b1101111000;  // alpha^120
            10'd 121: o_tuple = 10'b1011111001;  // alpha^121
            10'd 122: o_tuple = 10'b0111111011;  // alpha^122
            10'd 123: o_tuple = 10'b1111110110;  // alpha^123
            10'd 124: o_tuple = 10'b1111100101;  // alpha^124
            10'd 125: o_tuple = 10'b1111000011;  // alpha^125
            10'd 126: o_tuple = 10'b1110001111;  // alpha^126
            10'd 127: o_tuple = 10'b1100010111;  // alpha^127
            10'd 128: o_tuple = 10'b1000100111;  // alpha^128
            10'd 129: o_tuple = 10'b0001000111;  // alpha^129
            10'd 130: o_tuple = 10'b0010001110;  // alpha^130
            10'd 131: o_tuple = 10'b0100011100;  // alpha^131
            10'd 132: o_tuple = 10'b1000111000;  // alpha^132
            10'd 133: o_tuple = 10'b0001111001;  // alpha^133
            10'd 134: o_tuple = 10'b0011110010;  // alpha^134
            10'd 135: o_tuple = 10'b0111100100;  // alpha^135
            10'd 136: o_tuple = 10'b1111001000;  // alpha^136
            10'd 137: o_tuple = 10'b1110011001;  // alpha^137
            10'd 138: o_tuple = 10'b1100111011;  // alpha^138
            10'd 139: o_tuple = 10'b1001111111;  // alpha^139
            10'd 140: o_tuple = 10'b0011110111;  // alpha^140
            10'd 141: o_tuple = 10'b0111101110;  // alpha^141
            10'd 142: o_tuple = 10'b1111011100;  // alpha^142
            10'd 143: o_tuple = 10'b1110110001;  // alpha^143
            10'd 144: o_tuple = 10'b1101101011;  // alpha^144
            10'd 145: o_tuple = 10'b1011011111;  // alpha^145
            10'd 146: o_tuple = 10'b0110110111;  // alpha^146
            10'd 147: o_tuple = 10'b1101101110;  // alpha^147
            10'd 148: o_tuple = 10'b1011010101;  // alpha^148
            10'd 149: o_tuple = 10'b0110100011;  // alpha^149
            10'd 150: o_tuple = 10'b1101000110;  // alpha^150
            10'd 151: o_tuple = 10'b1010000101;  // alpha^151
            10'd 152: o_tuple = 10'b0100000011;  // alpha^152
            10'd 153: o_tuple = 10'b1000000110;  // alpha^153
            10'd 154: o_tuple = 10'b0000000101;  // alpha^154
            10'd 155: o_tuple = 10'b0000001010;  // alpha^155
            10'd 156: o_tuple = 10'b0000010100;  // alpha^156
            10'd 157: o_tuple = 10'b0000101000;  // alpha^157
            10'd 158: o_tuple = 10'b0001010000;  // alpha^158
            10'd 159: o_tuple = 10'b0010100000;  // alpha^159
            10'd 160: o_tuple = 10'b0101000000;  // alpha^160
            10'd 161: o_tuple = 10'b1010000000;  // alpha^161
            10'd 162: o_tuple = 10'b0100001001;  // alpha^162
            10'd 163: o_tuple = 10'b1000010010;  // alpha^163
            10'd 164: o_tuple = 10'b0000101101;  // alpha^164
            10'd 165: o_tuple = 10'b0001011010;  // alpha^165
            10'd 166: o_tuple = 10'b0010110100;  // alpha^166
            10'd 167: o_tuple = 10'b0101101000;  // alpha^167
            10'd 168: o_tuple = 10'b1011010000;  // alpha^168
            10'd 169: o_tuple = 10'b0110101001;  // alpha^169
            10'd 170: o_tuple = 10'b1101010010;  // alpha^170
            10'd 171: o_tuple = 10'b1010101101;  // alpha^171
            10'd 172: o_tuple = 10'b0101010011;  // alpha^172
            10'd 173: o_tuple = 10'b1010100110;  // alpha^173
            10'd 174: o_tuple = 10'b0101000101;  // alpha^174
            10'd 175: o_tuple = 10'b1010001010;  // alpha^175
            10'd 176: o_tuple = 10'b0100011101;  // alpha^176
            10'd 177: o_tuple = 10'b1000111010;  // alpha^177
            10'd 178: o_tuple = 10'b0001111101;  // alpha^178
            10'd 179: o_tuple = 10'b0011111010;  // alpha^179
            10'd 180: o_tuple = 10'b0111110100;  // alpha^180
            10'd 181: o_tuple = 10'b1111101000;  // alpha^181
            10'd 182: o_tuple = 10'b1111011001;  // alpha^182
            10'd 183: o_tuple = 10'b1110111011;  // alpha^183
            10'd 184: o_tuple = 10'b1101111111;  // alpha^184
            10'd 185: o_tuple = 10'b1011110111;  // alpha^185
            10'd 186: o_tuple = 10'b0111100111;  // alpha^186
            10'd 187: o_tuple = 10'b1111001110;  // alpha^187
            10'd 188: o_tuple = 10'b1110010101;  // alpha^188
            10'd 189: o_tuple = 10'b1100100011;  // alpha^189
            10'd 190: o_tuple = 10'b1001001111;  // alpha^190
            10'd 191: o_tuple = 10'b0010010111;  // alpha^191
            10'd 192: o_tuple = 10'b0100101110;  // alpha^192
            10'd 193: o_tuple = 10'b1001011100;  // alpha^193
            10'd 194: o_tuple = 10'b0010110001;  // alpha^194
            10'd 195: o_tuple = 10'b0101100010;  // alpha^195
            10'd 196: o_tuple = 10'b1011000100;  // alpha^196
            10'd 197: o_tuple = 10'b0110000001;  // alpha^197
            10'd 198: o_tuple = 10'b1100000010;  // alpha^198
            10'd 199: o_tuple = 10'b1000001101;  // alpha^199
            10'd 200: o_tuple = 10'b0000010011;  // alpha^200
            10'd 201: o_tuple = 10'b0000100110;  // alpha^201
            10'd 202: o_tuple = 10'b0001001100;  // alpha^202
            10'd 203: o_tuple = 10'b0010011000;  // alpha^203
            10'd 204: o_tuple = 10'b0100110000;  // alpha^204
            10'd 205: o_tuple = 10'b1001100000;  // alpha^205
            10'd 206: o_tuple = 10'b0011001001;  // alpha^206
            10'd 207: o_tuple = 10'b0110010010;  // alpha^207
            10'd 208: o_tuple = 10'b1100100100;  // alpha^208
            10'd 209: o_tuple = 10'b1001000001;  // alpha^209
            10'd 210: o_tuple = 10'b0010001011;  // alpha^210
            10'd 211: o_tuple = 10'b0100010110;  // alpha^211
            10'd 212: o_tuple = 10'b1000101100;  // alpha^212
            10'd 213: o_tuple = 10'b0001010001;  // alpha^213
            10'd 214: o_tuple = 10'b0010100010;  // alpha^214
            10'd 215: o_tuple = 10'b0101000100;  // alpha^215
            10'd 216: o_tuple = 10'b1010001000;  // alpha^216
            10'd 217: o_tuple = 10'b0100011001;  // alpha^217
            10'd 218: o_tuple = 10'b1000110010;  // alpha^218
            10'd 219: o_tuple = 10'b0001101101;  // alpha^219
            10'd 220: o_tuple = 10'b0011011010;  // alpha^220
            10'd 221: o_tuple = 10'b0110110100;  // alpha^221
            10'd 222: o_tuple = 10'b1101101000;  // alpha^222
            10'd 223: o_tuple = 10'b1011011001;  // alpha^223
            10'd 224: o_tuple = 10'b0110111011;  // alpha^224
            10'd 225: o_tuple = 10'b1101110110;  // alpha^225
            10'd 226: o_tuple = 10'b1011100101;  // alpha^226
            10'd 227: o_tuple = 10'b0111000011;  // alpha^227
            10'd 228: o_tuple = 10'b1110000110;  // alpha^228
            10'd 229: o_tuple = 10'b1100000101;  // alpha^229
            10'd 230: o_tuple = 10'b1000000011;  // alpha^230
            10'd 231: o_tuple = 10'b0000001111;  // alpha^231
            10'd 232: o_tuple = 10'b0000011110;  // alpha^232
            10'd 233: o_tuple = 10'b0000111100;  // alpha^233
            10'd 234: o_tuple = 10'b0001111000;  // alpha^234
            10'd 235: o_tuple = 10'b0011110000;  // alpha^235
            10'd 236: o_tuple = 10'b0111100000;  // alpha^236
            10'd 237: o_tuple = 10'b1111000000;  // alpha^237
            10'd 238: o_tuple = 10'b1110001001;  // alpha^238
            10'd 239: o_tuple = 10'b1100011011;  // alpha^239
            10'd 240: o_tuple = 10'b1000111111;  // alpha^240
            10'd 241: o_tuple = 10'b0001110111;  // alpha^241
            10'd 242: o_tuple = 10'b0011101110;  // alpha^242
            10'd 243: o_tuple = 10'b0111011100;  // alpha^243
            10'd 244: o_tuple = 10'b1110111000;  // alpha^244
            10'd 245: o_tuple = 10'b1101111001;  // alpha^245
            10'd 246: o_tuple = 10'b1011111011;  // alpha^246
            10'd 247: o_tuple = 10'b0111111111;  // alpha^247
            10'd 248: o_tuple = 10'b1111111110;  // alpha^248
            10'd 249: o_tuple = 10'b1111110101;  // alpha^249
            10'd 250: o_tuple = 10'b1111100011;  // alpha^250
            10'd 251: o_tuple = 10'b1111001111;  // alpha^251
            10'd 252: o_tuple = 10'b1110010111;  // alpha^252
            10'd 253: o_tuple = 10'b1100100111;  // alpha^253
            10'd 254: o_tuple = 10'b1001000111;  // alpha^254
            10'd 255: o_tuple = 10'b0010000111;  // alpha^255
            10'd 256: o_tuple = 10'b0100001110;  // alpha^256
            10'd 257: o_tuple = 10'b1000011100;  // alpha^257
            10'd 258: o_tuple = 10'b0000110001;  // alpha^258
            10'd 259: o_tuple = 10'b0001100010;  // alpha^259
            10'd 260: o_tuple = 10'b0011000100;  // alpha^260
            10'd 261: o_tuple = 10'b0110001000;  // alpha^261
            10'd 262: o_tuple = 10'b1100010000;  // alpha^262
            10'd 263: o_tuple = 10'b1000101001;  // alpha^263
            10'd 264: o_tuple = 10'b0001011011;  // alpha^264
            10'd 265: o_tuple = 10'b0010110110;  // alpha^265
            10'd 266: o_tuple = 10'b0101101100;  // alpha^266
            10'd 267: o_tuple = 10'b1011011000;  // alpha^267
            10'd 268: o_tuple = 10'b0110111001;  // alpha^268
            10'd 269: o_tuple = 10'b1101110010;  // alpha^269
            10'd 270: o_tuple = 10'b1011101101;  // alpha^270
            10'd 271: o_tuple = 10'b0111010011;  // alpha^271
            10'd 272: o_tuple = 10'b1110100110;  // alpha^272
            10'd 273: o_tuple = 10'b1101000101;  // alpha^273
            10'd 274: o_tuple = 10'b1010000011;  // alpha^274
            10'd 275: o_tuple = 10'b0100001111;  // alpha^275
            10'd 276: o_tuple = 10'b1000011110;  // alpha^276
            10'd 277: o_tuple = 10'b0000110101;  // alpha^277
            10'd 278: o_tuple = 10'b0001101010;  // alpha^278
            10'd 279: o_tuple = 10'b0011010100;  // alpha^279
            10'd 280: o_tuple = 10'b0110101000;  // alpha^280
            10'd 281: o_tuple = 10'b1101010000;  // alpha^281
            10'd 282: o_tuple = 10'b1010101001;  // alpha^282
            10'd 283: o_tuple = 10'b0101011011;  // alpha^283
            10'd 284: o_tuple = 10'b1010110110;  // alpha^284
            10'd 285: o_tuple = 10'b0101100101;  // alpha^285
            10'd 286: o_tuple = 10'b1011001010;  // alpha^286
            10'd 287: o_tuple = 10'b0110011101;  // alpha^287
            10'd 288: o_tuple = 10'b1100111010;  // alpha^288
            10'd 289: o_tuple = 10'b1001111101;  // alpha^289
            10'd 290: o_tuple = 10'b0011110011;  // alpha^290
            10'd 291: o_tuple = 10'b0111100110;  // alpha^291
            10'd 292: o_tuple = 10'b1111001100;  // alpha^292
            10'd 293: o_tuple = 10'b1110010001;  // alpha^293
            10'd 294: o_tuple = 10'b1100101011;  // alpha^294
            10'd 295: o_tuple = 10'b1001011111;  // alpha^295
            10'd 296: o_tuple = 10'b0010110111;  // alpha^296
            10'd 297: o_tuple = 10'b0101101110;  // alpha^297
            10'd 298: o_tuple = 10'b1011011100;  // alpha^298
            10'd 299: o_tuple = 10'b0110110001;  // alpha^299
            10'd 300: o_tuple = 10'b1101100010;  // alpha^300
            10'd 301: o_tuple = 10'b1011001101;  // alpha^301
            10'd 302: o_tuple = 10'b0110010011;  // alpha^302
            10'd 303: o_tuple = 10'b1100100110;  // alpha^303
            10'd 304: o_tuple = 10'b1001000101;  // alpha^304
            10'd 305: o_tuple = 10'b0010000011;  // alpha^305
            10'd 306: o_tuple = 10'b0100000110;  // alpha^306
            10'd 307: o_tuple = 10'b1000001100;  // alpha^307
            10'd 308: o_tuple = 10'b0000010001;  // alpha^308
            10'd 309: o_tuple = 10'b0000100010;  // alpha^309
            10'd 310: o_tuple = 10'b0001000100;  // alpha^310
            10'd 311: o_tuple = 10'b0010001000;  // alpha^311
            10'd 312: o_tuple = 10'b0100010000;  // alpha^312
            10'd 313: o_tuple = 10'b1000100000;  // alpha^313
            10'd 314: o_tuple = 10'b0001001001;  // alpha^314
            10'd 315: o_tuple = 10'b0010010010;  // alpha^315
            10'd 316: o_tuple = 10'b0100100100;  // alpha^316
            10'd 317: o_tuple = 10'b1001001000;  // alpha^317
            10'd 318: o_tuple = 10'b0010011001;  // alpha^318
            10'd 319: o_tuple = 10'b0100110010;  // alpha^319
            10'd 320: o_tuple = 10'b1001100100;  // alpha^320
            10'd 321: o_tuple = 10'b0011000001;  // alpha^321
            10'd 322: o_tuple = 10'b0110000010;  // alpha^322
            10'd 323: o_tuple = 10'b1100000100;  // alpha^323
            10'd 324: o_tuple = 10'b1000000001;  // alpha^324
            10'd 325: o_tuple = 10'b0000001011;  // alpha^325
            10'd 326: o_tuple = 10'b0000010110;  // alpha^326
            10'd 327: o_tuple = 10'b0000101100;  // alpha^327
            10'd 328: o_tuple = 10'b0001011000;  // alpha^328
            10'd 329: o_tuple = 10'b0010110000;  // alpha^329
            10'd 330: o_tuple = 10'b0101100000;  // alpha^330
            10'd 331: o_tuple = 10'b1011000000;  // alpha^331
            10'd 332: o_tuple = 10'b0110001001;  // alpha^332
            10'd 333: o_tuple = 10'b1100010010;  // alpha^333
            10'd 334: o_tuple = 10'b1000101101;  // alpha^334
            10'd 335: o_tuple = 10'b0001010011;  // alpha^335
            10'd 336: o_tuple = 10'b0010100110;  // alpha^336
            10'd 337: o_tuple = 10'b0101001100;  // alpha^337
            10'd 338: o_tuple = 10'b1010011000;  // alpha^338
            10'd 339: o_tuple = 10'b0100111001;  // alpha^339
            10'd 340: o_tuple = 10'b1001110010;  // alpha^340
            10'd 341: o_tuple = 10'b0011101101;  // alpha^341
            10'd 342: o_tuple = 10'b0111011010;  // alpha^342
            10'd 343: o_tuple = 10'b1110110100;  // alpha^343
            10'd 344: o_tuple = 10'b1101100001;  // alpha^344
            10'd 345: o_tuple = 10'b1011001011;  // alpha^345
            10'd 346: o_tuple = 10'b0110011111;  // alpha^346
            10'd 347: o_tuple = 10'b1100111110;  // alpha^347
            10'd 348: o_tuple = 10'b1001110101;  // alpha^348
            10'd 349: o_tuple = 10'b0011100011;  // alpha^349
            10'd 350: o_tuple = 10'b0111000110;  // alpha^350
            10'd 351: o_tuple = 10'b1110001100;  // alpha^351
            10'd 352: o_tuple = 10'b1100010001;  // alpha^352
            10'd 353: o_tuple = 10'b1000101011;  // alpha^353
            10'd 354: o_tuple = 10'b0001011111;  // alpha^354
            10'd 355: o_tuple = 10'b0010111110;  // alpha^355
            10'd 356: o_tuple = 10'b0101111100;  // alpha^356
            10'd 357: o_tuple = 10'b1011111000;  // alpha^357
            10'd 358: o_tuple = 10'b0111111001;  // alpha^358
            10'd 359: o_tuple = 10'b1111110010;  // alpha^359
            10'd 360: o_tuple = 10'b1111101101;  // alpha^360
            10'd 361: o_tuple = 10'b1111010011;  // alpha^361
            10'd 362: o_tuple = 10'b1110101111;  // alpha^362
            10'd 363: o_tuple = 10'b1101010111;  // alpha^363
            10'd 364: o_tuple = 10'b1010100111;  // alpha^364
            10'd 365: o_tuple = 10'b0101000111;  // alpha^365
            10'd 366: o_tuple = 10'b1010001110;  // alpha^366
            10'd 367: o_tuple = 10'b0100010101;  // alpha^367
            10'd 368: o_tuple = 10'b1000101010;  // alpha^368
            10'd 369: o_tuple = 10'b0001011101;  // alpha^369
            10'd 370: o_tuple = 10'b0010111010;  // alpha^370
            10'd 371: o_tuple = 10'b0101110100;  // alpha^371
            10'd 372: o_tuple = 10'b1011101000;  // alpha^372
            10'd 373: o_tuple = 10'b0111011001;  // alpha^373
            10'd 374: o_tuple = 10'b1110110010;  // alpha^374
            10'd 375: o_tuple = 10'b1101101101;  // alpha^375
            10'd 376: o_tuple = 10'b1011010011;  // alpha^376
            10'd 377: o_tuple = 10'b0110101111;  // alpha^377
            10'd 378: o_tuple = 10'b1101011110;  // alpha^378
            10'd 379: o_tuple = 10'b1010110101;  // alpha^379
            10'd 380: o_tuple = 10'b0101100011;  // alpha^380
            10'd 381: o_tuple = 10'b1011000110;  // alpha^381
            10'd 382: o_tuple = 10'b0110000101;  // alpha^382
            10'd 383: o_tuple = 10'b1100001010;  // alpha^383
            10'd 384: o_tuple = 10'b1000011101;  // alpha^384
            10'd 385: o_tuple = 10'b0000110011;  // alpha^385
            10'd 386: o_tuple = 10'b0001100110;  // alpha^386
            10'd 387: o_tuple = 10'b0011001100;  // alpha^387
            10'd 388: o_tuple = 10'b0110011000;  // alpha^388
            10'd 389: o_tuple = 10'b1100110000;  // alpha^389
            10'd 390: o_tuple = 10'b1001101001;  // alpha^390
            10'd 391: o_tuple = 10'b0011011011;  // alpha^391
            10'd 392: o_tuple = 10'b0110110110;  // alpha^392
            10'd 393: o_tuple = 10'b1101101100;  // alpha^393
            10'd 394: o_tuple = 10'b1011010001;  // alpha^394
            10'd 395: o_tuple = 10'b0110101011;  // alpha^395
            10'd 396: o_tuple = 10'b1101010110;  // alpha^396
            10'd 397: o_tuple = 10'b1010100101;  // alpha^397
            10'd 398: o_tuple = 10'b0101000011;  // alpha^398
            10'd 399: o_tuple = 10'b1010000110;  // alpha^399
            10'd 400: o_tuple = 10'b0100000101;  // alpha^400
            10'd 401: o_tuple = 10'b1000001010;  // alpha^401
            10'd 402: o_tuple = 10'b0000011101;  // alpha^402
            10'd 403: o_tuple = 10'b0000111010;  // alpha^403
            10'd 404: o_tuple = 10'b0001110100;  // alpha^404
            10'd 405: o_tuple = 10'b0011101000;  // alpha^405
            10'd 406: o_tuple = 10'b0111010000;  // alpha^406
            10'd 407: o_tuple = 10'b1110100000;  // alpha^407
            10'd 408: o_tuple = 10'b1101001001;  // alpha^408
            10'd 409: o_tuple = 10'b1010011011;  // alpha^409
            10'd 410: o_tuple = 10'b0100111111;  // alpha^410
            10'd 411: o_tuple = 10'b1001111110;  // alpha^411
            10'd 412: o_tuple = 10'b0011110101;  // alpha^412
            10'd 413: o_tuple = 10'b0111101010;  // alpha^413
            10'd 414: o_tuple = 10'b1111010100;  // alpha^414
            10'd 415: o_tuple = 10'b1110100001;  // alpha^415
            10'd 416: o_tuple = 10'b1101001011;  // alpha^416
            10'd 417: o_tuple = 10'b1010011111;  // alpha^417
            10'd 418: o_tuple = 10'b0100110111;  // alpha^418
            10'd 419: o_tuple = 10'b1001101110;  // alpha^419
            10'd 420: o_tuple = 10'b0011010101;  // alpha^420
            10'd 421: o_tuple = 10'b0110101010;  // alpha^421
            10'd 422: o_tuple = 10'b1101010100;  // alpha^422
            10'd 423: o_tuple = 10'b1010100001;  // alpha^423
            10'd 424: o_tuple = 10'b0101001011;  // alpha^424
            10'd 425: o_tuple = 10'b1010010110;  // alpha^425
            10'd 426: o_tuple = 10'b0100100101;  // alpha^426
            10'd 427: o_tuple = 10'b1001001010;  // alpha^427
            10'd 428: o_tuple = 10'b0010011101;  // alpha^428
            10'd 429: o_tuple = 10'b0100111010;  // alpha^429
            10'd 430: o_tuple = 10'b1001110100;  // alpha^430
            10'd 431: o_tuple = 10'b0011100001;  // alpha^431
            10'd 432: o_tuple = 10'b0111000010;  // alpha^432
            10'd 433: o_tuple = 10'b1110000100;  // alpha^433
            10'd 434: o_tuple = 10'b1100000001;  // alpha^434
            10'd 435: o_tuple = 10'b1000001011;  // alpha^435
            10'd 436: o_tuple = 10'b0000011111;  // alpha^436
            10'd 437: o_tuple = 10'b0000111110;  // alpha^437
            10'd 438: o_tuple = 10'b0001111100;  // alpha^438
            10'd 439: o_tuple = 10'b0011111000;  // alpha^439
            10'd 440: o_tuple = 10'b0111110000;  // alpha^440
            10'd 441: o_tuple = 10'b1111100000;  // alpha^441
            10'd 442: o_tuple = 10'b1111001001;  // alpha^442
            10'd 443: o_tuple = 10'b1110011011;  // alpha^443
            10'd 444: o_tuple = 10'b1100111111;  // alpha^444
            10'd 445: o_tuple = 10'b1001110111;  // alpha^445
            10'd 446: o_tuple = 10'b0011100111;  // alpha^446
            10'd 447: o_tuple = 10'b0111001110;  // alpha^447
            10'd 448: o_tuple = 10'b1110011100;  // alpha^448
            10'd 449: o_tuple = 10'b1100110001;  // alpha^449
            10'd 450: o_tuple = 10'b1001101011;  // alpha^450
            10'd 451: o_tuple = 10'b0011011111;  // alpha^451
            10'd 452: o_tuple = 10'b0110111110;  // alpha^452
            10'd 453: o_tuple = 10'b1101111100;  // alpha^453
            10'd 454: o_tuple = 10'b1011110001;  // alpha^454
            10'd 455: o_tuple = 10'b0111101011;  // alpha^455
            10'd 456: o_tuple = 10'b1111010110;  // alpha^456
            10'd 457: o_tuple = 10'b1110100101;  // alpha^457
            10'd 458: o_tuple = 10'b1101000011;  // alpha^458
            10'd 459: o_tuple = 10'b1010001111;  // alpha^459
            10'd 460: o_tuple = 10'b0100010111;  // alpha^460
            10'd 461: o_tuple = 10'b1000101110;  // alpha^461
            10'd 462: o_tuple = 10'b0001010101;  // alpha^462
            10'd 463: o_tuple = 10'b0010101010;  // alpha^463
            10'd 464: o_tuple = 10'b0101010100;  // alpha^464
            10'd 465: o_tuple = 10'b1010101000;  // alpha^465
            10'd 466: o_tuple = 10'b0101011001;  // alpha^466
            10'd 467: o_tuple = 10'b1010110010;  // alpha^467
            10'd 468: o_tuple = 10'b0101101101;  // alpha^468
            10'd 469: o_tuple = 10'b1011011010;  // alpha^469
            10'd 470: o_tuple = 10'b0110111101;  // alpha^470
            10'd 471: o_tuple = 10'b1101111010;  // alpha^471
            10'd 472: o_tuple = 10'b1011111101;  // alpha^472
            10'd 473: o_tuple = 10'b0111110011;  // alpha^473
            10'd 474: o_tuple = 10'b1111100110;  // alpha^474
            10'd 475: o_tuple = 10'b1111000101;  // alpha^475
            10'd 476: o_tuple = 10'b1110000011;  // alpha^476
            10'd 477: o_tuple = 10'b1100001111;  // alpha^477
            10'd 478: o_tuple = 10'b1000010111;  // alpha^478
            10'd 479: o_tuple = 10'b0000100111;  // alpha^479
            10'd 480: o_tuple = 10'b0001001110;  // alpha^480
            10'd 481: o_tuple = 10'b0010011100;  // alpha^481
            10'd 482: o_tuple = 10'b0100111000;  // alpha^482
            10'd 483: o_tuple = 10'b1001110000;  // alpha^483
            10'd 484: o_tuple = 10'b0011101001;  // alpha^484
            10'd 485: o_tuple = 10'b0111010010;  // alpha^485
            10'd 486: o_tuple = 10'b1110100100;  // alpha^486
            10'd 487: o_tuple = 10'b1101000001;  // alpha^487
            10'd 488: o_tuple = 10'b1010001011;  // alpha^488
            10'd 489: o_tuple = 10'b0100011111;  // alpha^489
            10'd 490: o_tuple = 10'b1000111110;  // alpha^490
            10'd 491: o_tuple = 10'b0001110101;  // alpha^491
            10'd 492: o_tuple = 10'b0011101010;  // alpha^492
            10'd 493: o_tuple = 10'b0111010100;  // alpha^493
            10'd 494: o_tuple = 10'b1110101000;  // alpha^494
            10'd 495: o_tuple = 10'b1101011001;  // alpha^495
            10'd 496: o_tuple = 10'b1010111011;  // alpha^496
            10'd 497: o_tuple = 10'b0101111111;  // alpha^497
            10'd 498: o_tuple = 10'b1011111110;  // alpha^498
            10'd 499: o_tuple = 10'b0111110101;  // alpha^499
            10'd 500: o_tuple = 10'b1111101010;  // alpha^500
            10'd 501: o_tuple = 10'b1111011101;  // alpha^501
            10'd 502: o_tuple = 10'b1110110011;  // alpha^502
            10'd 503: o_tuple = 10'b1101101111;  // alpha^503
            10'd 504: o_tuple = 10'b1011010111;  // alpha^504
            10'd 505: o_tuple = 10'b0110100111;  // alpha^505
            10'd 506: o_tuple = 10'b1101001110;  // alpha^506
            10'd 507: o_tuple = 10'b1010010101;  // alpha^507
            10'd 508: o_tuple = 10'b0100100011;  // alpha^508
            10'd 509: o_tuple = 10'b1001000110;  // alpha^509
            10'd 510: o_tuple = 10'b0010000101;  // alpha^510
            10'd 511: o_tuple = 10'b0100001010;  // alpha^511
            10'd 512: o_tuple = 10'b1000010100;  // alpha^512
            10'd 513: o_tuple = 10'b0000100001;  // alpha^513
            10'd 514: o_tuple = 10'b0001000010;  // alpha^514
            10'd 515: o_tuple = 10'b0010000100;  // alpha^515
            10'd 516: o_tuple = 10'b0100001000;  // alpha^516
            10'd 517: o_tuple = 10'b1000010000;  // alpha^517
            10'd 518: o_tuple = 10'b0000101001;  // alpha^518
            10'd 519: o_tuple = 10'b0001010010;  // alpha^519
            10'd 520: o_tuple = 10'b0010100100;  // alpha^520
            10'd 521: o_tuple = 10'b0101001000;  // alpha^521
            10'd 522: o_tuple = 10'b1010010000;  // alpha^522
            10'd 523: o_tuple = 10'b0100101001;  // alpha^523
            10'd 524: o_tuple = 10'b1001010010;  // alpha^524
            10'd 525: o_tuple = 10'b0010101101;  // alpha^525
            10'd 526: o_tuple = 10'b0101011010;  // alpha^526
            10'd 527: o_tuple = 10'b1010110100;  // alpha^527
            10'd 528: o_tuple = 10'b0101100001;  // alpha^528
            10'd 529: o_tuple = 10'b1011000010;  // alpha^529
            10'd 530: o_tuple = 10'b0110001101;  // alpha^530
            10'd 531: o_tuple = 10'b1100011010;  // alpha^531
            10'd 532: o_tuple = 10'b1000111101;  // alpha^532
            10'd 533: o_tuple = 10'b0001110011;  // alpha^533
            10'd 534: o_tuple = 10'b0011100110;  // alpha^534
            10'd 535: o_tuple = 10'b0111001100;  // alpha^535
            10'd 536: o_tuple = 10'b1110011000;  // alpha^536
            10'd 537: o_tuple = 10'b1100111001;  // alpha^537
            10'd 538: o_tuple = 10'b1001111011;  // alpha^538
            10'd 539: o_tuple = 10'b0011111111;  // alpha^539
            10'd 540: o_tuple = 10'b0111111110;  // alpha^540
            10'd 541: o_tuple = 10'b1111111100;  // alpha^541
            10'd 542: o_tuple = 10'b1111110001;  // alpha^542
            10'd 543: o_tuple = 10'b1111101011;  // alpha^543
            10'd 544: o_tuple = 10'b1111011111;  // alpha^544
            10'd 545: o_tuple = 10'b1110110111;  // alpha^545
            10'd 546: o_tuple = 10'b1101100111;  // alpha^546
            10'd 547: o_tuple = 10'b1011000111;  // alpha^547
            10'd 548: o_tuple = 10'b0110000111;  // alpha^548
            10'd 549: o_tuple = 10'b1100001110;  // alpha^549
            10'd 550: o_tuple = 10'b1000010101;  // alpha^550
            10'd 551: o_tuple = 10'b0000100011;  // alpha^551
            10'd 552: o_tuple = 10'b0001000110;  // alpha^552
            10'd 553: o_tuple = 10'b0010001100;  // alpha^553
            10'd 554: o_tuple = 10'b0100011000;  // alpha^554
            10'd 555: o_tuple = 10'b1000110000;  // alpha^555
            10'd 556: o_tuple = 10'b0001101001;  // alpha^556
            10'd 557: o_tuple = 10'b0011010010;  // alpha^557
            10'd 558: o_tuple = 10'b0110100100;  // alpha^558
            10'd 559: o_tuple = 10'b1101001000;  // alpha^559
            10'd 560: o_tuple = 10'b1010011001;  // alpha^560
            10'd 561: o_tuple = 10'b0100111011;  // alpha^561
            10'd 562: o_tuple = 10'b1001110110;  // alpha^562
            10'd 563: o_tuple = 10'b0011100101;  // alpha^563
            10'd 564: o_tuple = 10'b0111001010;  // alpha^564
            10'd 565: o_tuple = 10'b1110010100;  // alpha^565
            10'd 566: o_tuple = 10'b1100100001;  // alpha^566
            10'd 567: o_tuple = 10'b1001001011;  // alpha^567
            10'd 568: o_tuple = 10'b0010011111;  // alpha^568
            10'd 569: o_tuple = 10'b0100111110;  // alpha^569
            10'd 570: o_tuple = 10'b1001111100;  // alpha^570
            10'd 571: o_tuple = 10'b0011110001;  // alpha^571
            10'd 572: o_tuple = 10'b0111100010;  // alpha^572
            10'd 573: o_tuple = 10'b1111000100;  // alpha^573
            10'd 574: o_tuple = 10'b1110000001;  // alpha^574
            10'd 575: o_tuple = 10'b1100001011;  // alpha^575
            10'd 576: o_tuple = 10'b1000011111;  // alpha^576
            10'd 577: o_tuple = 10'b0000110111;  // alpha^577
            10'd 578: o_tuple = 10'b0001101110;  // alpha^578
            10'd 579: o_tuple = 10'b0011011100;  // alpha^579
            10'd 580: o_tuple = 10'b0110111000;  // alpha^580
            10'd 581: o_tuple = 10'b1101110000;  // alpha^581
            10'd 582: o_tuple = 10'b1011101001;  // alpha^582
            10'd 583: o_tuple = 10'b0111011011;  // alpha^583
            10'd 584: o_tuple = 10'b1110110110;  // alpha^584
            10'd 585: o_tuple = 10'b1101100101;  // alpha^585
            10'd 586: o_tuple = 10'b1011000011;  // alpha^586
            10'd 587: o_tuple = 10'b0110001111;  // alpha^587
            10'd 588: o_tuple = 10'b1100011110;  // alpha^588
            10'd 589: o_tuple = 10'b1000110101;  // alpha^589
            10'd 590: o_tuple = 10'b0001100011;  // alpha^590
            10'd 591: o_tuple = 10'b0011000110;  // alpha^591
            10'd 592: o_tuple = 10'b0110001100;  // alpha^592
            10'd 593: o_tuple = 10'b1100011000;  // alpha^593
            10'd 594: o_tuple = 10'b1000111001;  // alpha^594
            10'd 595: o_tuple = 10'b0001111011;  // alpha^595
            10'd 596: o_tuple = 10'b0011110110;  // alpha^596
            10'd 597: o_tuple = 10'b0111101100;  // alpha^597
            10'd 598: o_tuple = 10'b1111011000;  // alpha^598
            10'd 599: o_tuple = 10'b1110111001;  // alpha^599
            10'd 600: o_tuple = 10'b1101111011;  // alpha^600
            10'd 601: o_tuple = 10'b1011111111;  // alpha^601
            10'd 602: o_tuple = 10'b0111110111;  // alpha^602
            10'd 603: o_tuple = 10'b1111101110;  // alpha^603
            10'd 604: o_tuple = 10'b1111010101;  // alpha^604
            10'd 605: o_tuple = 10'b1110100011;  // alpha^605
            10'd 606: o_tuple = 10'b1101001111;  // alpha^606
            10'd 607: o_tuple = 10'b1010010111;  // alpha^607
            10'd 608: o_tuple = 10'b0100100111;  // alpha^608
            10'd 609: o_tuple = 10'b1001001110;  // alpha^609
            10'd 610: o_tuple = 10'b0010010101;  // alpha^610
            10'd 611: o_tuple = 10'b0100101010;  // alpha^611
            10'd 612: o_tuple = 10'b1001010100;  // alpha^612
            10'd 613: o_tuple = 10'b0010100001;  // alpha^613
            10'd 614: o_tuple = 10'b0101000010;  // alpha^614
            10'd 615: o_tuple = 10'b1010000100;  // alpha^615
            10'd 616: o_tuple = 10'b0100000001;  // alpha^616
            10'd 617: o_tuple = 10'b1000000010;  // alpha^617
            10'd 618: o_tuple = 10'b0000001101;  // alpha^618
            10'd 619: o_tuple = 10'b0000011010;  // alpha^619
            10'd 620: o_tuple = 10'b0000110100;  // alpha^620
            10'd 621: o_tuple = 10'b0001101000;  // alpha^621
            10'd 622: o_tuple = 10'b0011010000;  // alpha^622
            10'd 623: o_tuple = 10'b0110100000;  // alpha^623
            10'd 624: o_tuple = 10'b1101000000;  // alpha^624
            10'd 625: o_tuple = 10'b1010001001;  // alpha^625
            10'd 626: o_tuple = 10'b0100011011;  // alpha^626
            10'd 627: o_tuple = 10'b1000110110;  // alpha^627
            10'd 628: o_tuple = 10'b0001100101;  // alpha^628
            10'd 629: o_tuple = 10'b0011001010;  // alpha^629
            10'd 630: o_tuple = 10'b0110010100;  // alpha^630
            10'd 631: o_tuple = 10'b1100101000;  // alpha^631
            10'd 632: o_tuple = 10'b1001011001;  // alpha^632
            10'd 633: o_tuple = 10'b0010111011;  // alpha^633
            10'd 634: o_tuple = 10'b0101110110;  // alpha^634
            10'd 635: o_tuple = 10'b1011101100;  // alpha^635
            10'd 636: o_tuple = 10'b0111010001;  // alpha^636
            10'd 637: o_tuple = 10'b1110100010;  // alpha^637
            10'd 638: o_tuple = 10'b1101001101;  // alpha^638
            10'd 639: o_tuple = 10'b1010010011;  // alpha^639
            10'd 640: o_tuple = 10'b0100101111;  // alpha^640
            10'd 641: o_tuple = 10'b1001011110;  // alpha^641
            10'd 642: o_tuple = 10'b0010110101;  // alpha^642
            10'd 643: o_tuple = 10'b0101101010;  // alpha^643
            10'd 644: o_tuple = 10'b1011010100;  // alpha^644
            10'd 645: o_tuple = 10'b0110100001;  // alpha^645
            10'd 646: o_tuple = 10'b1101000010;  // alpha^646
            10'd 647: o_tuple = 10'b1010001101;  // alpha^647
            10'd 648: o_tuple = 10'b0100010011;  // alpha^648
            10'd 649: o_tuple = 10'b1000100110;  // alpha^649
            10'd 650: o_tuple = 10'b0001000101;  // alpha^650
            10'd 651: o_tuple = 10'b0010001010;  // alpha^651
            10'd 652: o_tuple = 10'b0100010100;  // alpha^652
            10'd 653: o_tuple = 10'b1000101000;  // alpha^653
            10'd 654: o_tuple = 10'b0001011001;  // alpha^654
            10'd 655: o_tuple = 10'b0010110010;  // alpha^655
            10'd 656: o_tuple = 10'b0101100100;  // alpha^656
            10'd 657: o_tuple = 10'b1011001000;  // alpha^657
            10'd 658: o_tuple = 10'b0110011001;  // alpha^658
            10'd 659: o_tuple = 10'b1100110010;  // alpha^659
            10'd 660: o_tuple = 10'b1001101101;  // alpha^660
            10'd 661: o_tuple = 10'b0011010011;  // alpha^661
            10'd 662: o_tuple = 10'b0110100110;  // alpha^662
            10'd 663: o_tuple = 10'b1101001100;  // alpha^663
            10'd 664: o_tuple = 10'b1010010001;  // alpha^664
            10'd 665: o_tuple = 10'b0100101011;  // alpha^665
            10'd 666: o_tuple = 10'b1001010110;  // alpha^666
            10'd 667: o_tuple = 10'b0010100101;  // alpha^667
            10'd 668: o_tuple = 10'b0101001010;  // alpha^668
            10'd 669: o_tuple = 10'b1010010100;  // alpha^669
            10'd 670: o_tuple = 10'b0100100001;  // alpha^670
            10'd 671: o_tuple = 10'b1001000010;  // alpha^671
            10'd 672: o_tuple = 10'b0010001101;  // alpha^672
            10'd 673: o_tuple = 10'b0100011010;  // alpha^673
            10'd 674: o_tuple = 10'b1000110100;  // alpha^674
            10'd 675: o_tuple = 10'b0001100001;  // alpha^675
            10'd 676: o_tuple = 10'b0011000010;  // alpha^676
            10'd 677: o_tuple = 10'b0110000100;  // alpha^677
            10'd 678: o_tuple = 10'b1100001000;  // alpha^678
            10'd 679: o_tuple = 10'b1000011001;  // alpha^679
            10'd 680: o_tuple = 10'b0000111011;  // alpha^680
            10'd 681: o_tuple = 10'b0001110110;  // alpha^681
            10'd 682: o_tuple = 10'b0011101100;  // alpha^682
            10'd 683: o_tuple = 10'b0111011000;  // alpha^683
            10'd 684: o_tuple = 10'b1110110000;  // alpha^684
            10'd 685: o_tuple = 10'b1101101001;  // alpha^685
            10'd 686: o_tuple = 10'b1011011011;  // alpha^686
            10'd 687: o_tuple = 10'b0110111111;  // alpha^687
            10'd 688: o_tuple = 10'b1101111110;  // alpha^688
            10'd 689: o_tuple = 10'b1011110101;  // alpha^689
            10'd 690: o_tuple = 10'b0111100011;  // alpha^690
            10'd 691: o_tuple = 10'b1111000110;  // alpha^691
            10'd 692: o_tuple = 10'b1110000101;  // alpha^692
            10'd 693: o_tuple = 10'b1100000011;  // alpha^693
            10'd 694: o_tuple = 10'b1000001111;  // alpha^694
            10'd 695: o_tuple = 10'b0000010111;  // alpha^695
            10'd 696: o_tuple = 10'b0000101110;  // alpha^696
            10'd 697: o_tuple = 10'b0001011100;  // alpha^697
            10'd 698: o_tuple = 10'b0010111000;  // alpha^698
            10'd 699: o_tuple = 10'b0101110000;  // alpha^699
            10'd 700: o_tuple = 10'b1011100000;  // alpha^700
            10'd 701: o_tuple = 10'b0111001001;  // alpha^701
            10'd 702: o_tuple = 10'b1110010010;  // alpha^702
            10'd 703: o_tuple = 10'b1100101101;  // alpha^703
            10'd 704: o_tuple = 10'b1001010011;  // alpha^704
            10'd 705: o_tuple = 10'b0010101111;  // alpha^705
            10'd 706: o_tuple = 10'b0101011110;  // alpha^706
            10'd 707: o_tuple = 10'b1010111100;  // alpha^707
            10'd 708: o_tuple = 10'b0101110001;  // alpha^708
            10'd 709: o_tuple = 10'b1011100010;  // alpha^709
            10'd 710: o_tuple = 10'b0111001101;  // alpha^710
            10'd 711: o_tuple = 10'b1110011010;  // alpha^711
            10'd 712: o_tuple = 10'b1100111101;  // alpha^712
            10'd 713: o_tuple = 10'b1001110011;  // alpha^713
            10'd 714: o_tuple = 10'b0011101111;  // alpha^714
            10'd 715: o_tuple = 10'b0111011110;  // alpha^715
            10'd 716: o_tuple = 10'b1110111100;  // alpha^716
            10'd 717: o_tuple = 10'b1101110001;  // alpha^717
            10'd 718: o_tuple = 10'b1011101011;  // alpha^718
            10'd 719: o_tuple = 10'b0111011111;  // alpha^719
            10'd 720: o_tuple = 10'b1110111110;  // alpha^720
            10'd 721: o_tuple = 10'b1101110101;  // alpha^721
            10'd 722: o_tuple = 10'b1011100011;  // alpha^722
            10'd 723: o_tuple = 10'b0111001111;  // alpha^723
            10'd 724: o_tuple = 10'b1110011110;  // alpha^724
            10'd 725: o_tuple = 10'b1100110101;  // alpha^725
            10'd 726: o_tuple = 10'b1001100011;  // alpha^726
            10'd 727: o_tuple = 10'b0011001111;  // alpha^727
            10'd 728: o_tuple = 10'b0110011110;  // alpha^728
            10'd 729: o_tuple = 10'b1100111100;  // alpha^729
            10'd 730: o_tuple = 10'b1001110001;  // alpha^730
            10'd 731: o_tuple = 10'b0011101011;  // alpha^731
            10'd 732: o_tuple = 10'b0111010110;  // alpha^732
            10'd 733: o_tuple = 10'b1110101100;  // alpha^733
            10'd 734: o_tuple = 10'b1101010001;  // alpha^734
            10'd 735: o_tuple = 10'b1010101011;  // alpha^735
            10'd 736: o_tuple = 10'b0101011111;  // alpha^736
            10'd 737: o_tuple = 10'b1010111110;  // alpha^737
            10'd 738: o_tuple = 10'b0101110101;  // alpha^738
            10'd 739: o_tuple = 10'b1011101010;  // alpha^739
            10'd 740: o_tuple = 10'b0111011101;  // alpha^740
            10'd 741: o_tuple = 10'b1110111010;  // alpha^741
            10'd 742: o_tuple = 10'b1101111101;  // alpha^742
            10'd 743: o_tuple = 10'b1011110011;  // alpha^743
            10'd 744: o_tuple = 10'b0111101111;  // alpha^744
            10'd 745: o_tuple = 10'b1111011110;  // alpha^745
            10'd 746: o_tuple = 10'b1110110101;  // alpha^746
            10'd 747: o_tuple = 10'b1101100011;  // alpha^747
            10'd 748: o_tuple = 10'b1011001111;  // alpha^748
            10'd 749: o_tuple = 10'b0110010111;  // alpha^749
            10'd 750: o_tuple = 10'b1100101110;  // alpha^750
            10'd 751: o_tuple = 10'b1001010101;  // alpha^751
            10'd 752: o_tuple = 10'b0010100011;  // alpha^752
            10'd 753: o_tuple = 10'b0101000110;  // alpha^753
            10'd 754: o_tuple = 10'b1010001100;  // alpha^754
            10'd 755: o_tuple = 10'b0100010001;  // alpha^755
            10'd 756: o_tuple = 10'b1000100010;  // alpha^756
            10'd 757: o_tuple = 10'b0001001101;  // alpha^757
            10'd 758: o_tuple = 10'b0010011010;  // alpha^758
            10'd 759: o_tuple = 10'b0100110100;  // alpha^759
            10'd 760: o_tuple = 10'b1001101000;  // alpha^760
            10'd 761: o_tuple = 10'b0011011001;  // alpha^761
            10'd 762: o_tuple = 10'b0110110010;  // alpha^762
            10'd 763: o_tuple = 10'b1101100100;  // alpha^763
            10'd 764: o_tuple = 10'b1011000001;  // alpha^764
            10'd 765: o_tuple = 10'b0110001011;  // alpha^765
            10'd 766: o_tuple = 10'b1100010110;  // alpha^766
            10'd 767: o_tuple = 10'b1000100101;  // alpha^767
            10'd 768: o_tuple = 10'b0001000011;  // alpha^768
            10'd 769: o_tuple = 10'b0010000110;  // alpha^769
            10'd 770: o_tuple = 10'b0100001100;  // alpha^770
            10'd 771: o_tuple = 10'b1000011000;  // alpha^771
            10'd 772: o_tuple = 10'b0000111001;  // alpha^772
            10'd 773: o_tuple = 10'b0001110010;  // alpha^773
            10'd 774: o_tuple = 10'b0011100100;  // alpha^774
            10'd 775: o_tuple = 10'b0111001000;  // alpha^775
            10'd 776: o_tuple = 10'b1110010000;  // alpha^776
            10'd 777: o_tuple = 10'b1100101001;  // alpha^777
            10'd 778: o_tuple = 10'b1001011011;  // alpha^778
            10'd 779: o_tuple = 10'b0010111111;  // alpha^779
            10'd 780: o_tuple = 10'b0101111110;  // alpha^780
            10'd 781: o_tuple = 10'b1011111100;  // alpha^781
            10'd 782: o_tuple = 10'b0111110001;  // alpha^782
            10'd 783: o_tuple = 10'b1111100010;  // alpha^783
            10'd 784: o_tuple = 10'b1111001101;  // alpha^784
            10'd 785: o_tuple = 10'b1110010011;  // alpha^785
            10'd 786: o_tuple = 10'b1100101111;  // alpha^786
            10'd 787: o_tuple = 10'b1001010111;  // alpha^787
            10'd 788: o_tuple = 10'b0010100111;  // alpha^788
            10'd 789: o_tuple = 10'b0101001110;  // alpha^789
            10'd 790: o_tuple = 10'b1010011100;  // alpha^790
            10'd 791: o_tuple = 10'b0100110001;  // alpha^791
            10'd 792: o_tuple = 10'b1001100010;  // alpha^792
            10'd 793: o_tuple = 10'b0011001101;  // alpha^793
            10'd 794: o_tuple = 10'b0110011010;  // alpha^794
            10'd 795: o_tuple = 10'b1100110100;  // alpha^795
            10'd 796: o_tuple = 10'b1001100001;  // alpha^796
            10'd 797: o_tuple = 10'b0011001011;  // alpha^797
            10'd 798: o_tuple = 10'b0110010110;  // alpha^798
            10'd 799: o_tuple = 10'b1100101100;  // alpha^799
            10'd 800: o_tuple = 10'b1001010001;  // alpha^800
            10'd 801: o_tuple = 10'b0010101011;  // alpha^801
            10'd 802: o_tuple = 10'b0101010110;  // alpha^802
            10'd 803: o_tuple = 10'b1010101100;  // alpha^803
            10'd 804: o_tuple = 10'b0101010001;  // alpha^804
            10'd 805: o_tuple = 10'b1010100010;  // alpha^805
            10'd 806: o_tuple = 10'b0101001101;  // alpha^806
            10'd 807: o_tuple = 10'b1010011010;  // alpha^807
            10'd 808: o_tuple = 10'b0100111101;  // alpha^808
            10'd 809: o_tuple = 10'b1001111010;  // alpha^809
            10'd 810: o_tuple = 10'b0011111101;  // alpha^810
            10'd 811: o_tuple = 10'b0111111010;  // alpha^811
            10'd 812: o_tuple = 10'b1111110100;  // alpha^812
            10'd 813: o_tuple = 10'b1111100001;  // alpha^813
            10'd 814: o_tuple = 10'b1111001011;  // alpha^814
            10'd 815: o_tuple = 10'b1110011111;  // alpha^815
            10'd 816: o_tuple = 10'b1100110111;  // alpha^816
            10'd 817: o_tuple = 10'b1001100111;  // alpha^817
            10'd 818: o_tuple = 10'b0011000111;  // alpha^818
            10'd 819: o_tuple = 10'b0110001110;  // alpha^819
            10'd 820: o_tuple = 10'b1100011100;  // alpha^820
            10'd 821: o_tuple = 10'b1000110001;  // alpha^821
            10'd 822: o_tuple = 10'b0001101011;  // alpha^822
            10'd 823: o_tuple = 10'b0011010110;  // alpha^823
            10'd 824: o_tuple = 10'b0110101100;  // alpha^824
            10'd 825: o_tuple = 10'b1101011000;  // alpha^825
            10'd 826: o_tuple = 10'b1010111001;  // alpha^826
            10'd 827: o_tuple = 10'b0101111011;  // alpha^827
            10'd 828: o_tuple = 10'b1011110110;  // alpha^828
            10'd 829: o_tuple = 10'b0111100101;  // alpha^829
            10'd 830: o_tuple = 10'b1111001010;  // alpha^830
            10'd 831: o_tuple = 10'b1110011101;  // alpha^831
            10'd 832: o_tuple = 10'b1100110011;  // alpha^832
            10'd 833: o_tuple = 10'b1001101111;  // alpha^833
            10'd 834: o_tuple = 10'b0011010111;  // alpha^834
            10'd 835: o_tuple = 10'b0110101110;  // alpha^835
            10'd 836: o_tuple = 10'b1101011100;  // alpha^836
            10'd 837: o_tuple = 10'b1010110001;  // alpha^837
            10'd 838: o_tuple = 10'b0101101011;  // alpha^838
            10'd 839: o_tuple = 10'b1011010110;  // alpha^839
            10'd 840: o_tuple = 10'b0110100101;  // alpha^840
            10'd 841: o_tuple = 10'b1101001010;  // alpha^841
            10'd 842: o_tuple = 10'b1010011101;  // alpha^842
            10'd 843: o_tuple = 10'b0100110011;  // alpha^843
            10'd 844: o_tuple = 10'b1001100110;  // alpha^844
            10'd 845: o_tuple = 10'b0011000101;  // alpha^845
            10'd 846: o_tuple = 10'b0110001010;  // alpha^846
            10'd 847: o_tuple = 10'b1100010100;  // alpha^847
            10'd 848: o_tuple = 10'b1000100001;  // alpha^848
            10'd 849: o_tuple = 10'b0001001011;  // alpha^849
            10'd 850: o_tuple = 10'b0010010110;  // alpha^850
            10'd 851: o_tuple = 10'b0100101100;  // alpha^851
            10'd 852: o_tuple = 10'b1001011000;  // alpha^852
            10'd 853: o_tuple = 10'b0010111001;  // alpha^853
            10'd 854: o_tuple = 10'b0101110010;  // alpha^854
            10'd 855: o_tuple = 10'b1011100100;  // alpha^855
            10'd 856: o_tuple = 10'b0111000001;  // alpha^856
            10'd 857: o_tuple = 10'b1110000010;  // alpha^857
            10'd 858: o_tuple = 10'b1100001101;  // alpha^858
            10'd 859: o_tuple = 10'b1000010011;  // alpha^859
            10'd 860: o_tuple = 10'b0000101111;  // alpha^860
            10'd 861: o_tuple = 10'b0001011110;  // alpha^861
            10'd 862: o_tuple = 10'b0010111100;  // alpha^862
            10'd 863: o_tuple = 10'b0101111000;  // alpha^863
            10'd 864: o_tuple = 10'b1011110000;  // alpha^864
            10'd 865: o_tuple = 10'b0111101001;  // alpha^865
            10'd 866: o_tuple = 10'b1111010010;  // alpha^866
            10'd 867: o_tuple = 10'b1110101101;  // alpha^867
            10'd 868: o_tuple = 10'b1101010011;  // alpha^868
            10'd 869: o_tuple = 10'b1010101111;  // alpha^869
            10'd 870: o_tuple = 10'b0101010111;  // alpha^870
            10'd 871: o_tuple = 10'b1010101110;  // alpha^871
            10'd 872: o_tuple = 10'b0101010101;  // alpha^872
            10'd 873: o_tuple = 10'b1010101010;  // alpha^873
            10'd 874: o_tuple = 10'b0101011101;  // alpha^874
            10'd 875: o_tuple = 10'b1010111010;  // alpha^875
            10'd 876: o_tuple = 10'b0101111101;  // alpha^876
            10'd 877: o_tuple = 10'b1011111010;  // alpha^877
            10'd 878: o_tuple = 10'b0111111101;  // alpha^878
            10'd 879: o_tuple = 10'b1111111010;  // alpha^879
            10'd 880: o_tuple = 10'b1111111101;  // alpha^880
            10'd 881: o_tuple = 10'b1111110011;  // alpha^881
            10'd 882: o_tuple = 10'b1111101111;  // alpha^882
            10'd 883: o_tuple = 10'b1111010111;  // alpha^883
            10'd 884: o_tuple = 10'b1110100111;  // alpha^884
            10'd 885: o_tuple = 10'b1101000111;  // alpha^885
            10'd 886: o_tuple = 10'b1010000111;  // alpha^886
            10'd 887: o_tuple = 10'b0100000111;  // alpha^887
            10'd 888: o_tuple = 10'b1000001110;  // alpha^888
            10'd 889: o_tuple = 10'b0000010101;  // alpha^889
            10'd 890: o_tuple = 10'b0000101010;  // alpha^890
            10'd 891: o_tuple = 10'b0001010100;  // alpha^891
            10'd 892: o_tuple = 10'b0010101000;  // alpha^892
            10'd 893: o_tuple = 10'b0101010000;  // alpha^893
            10'd 894: o_tuple = 10'b1010100000;  // alpha^894
            10'd 895: o_tuple = 10'b0101001001;  // alpha^895
            10'd 896: o_tuple = 10'b1010010010;  // alpha^896
            10'd 897: o_tuple = 10'b0100101101;  // alpha^897
            10'd 898: o_tuple = 10'b1001011010;  // alpha^898
            10'd 899: o_tuple = 10'b0010111101;  // alpha^899
            10'd 900: o_tuple = 10'b0101111010;  // alpha^900
            10'd 901: o_tuple = 10'b1011110100;  // alpha^901
            10'd 902: o_tuple = 10'b0111100001;  // alpha^902
            10'd 903: o_tuple = 10'b1111000010;  // alpha^903
            10'd 904: o_tuple = 10'b1110001101;  // alpha^904
            10'd 905: o_tuple = 10'b1100010011;  // alpha^905
            10'd 906: o_tuple = 10'b1000101111;  // alpha^906
            10'd 907: o_tuple = 10'b0001010111;  // alpha^907
            10'd 908: o_tuple = 10'b0010101110;  // alpha^908
            10'd 909: o_tuple = 10'b0101011100;  // alpha^909
            10'd 910: o_tuple = 10'b1010111000;  // alpha^910
            10'd 911: o_tuple = 10'b0101111001;  // alpha^911
            10'd 912: o_tuple = 10'b1011110010;  // alpha^912
            10'd 913: o_tuple = 10'b0111101101;  // alpha^913
            10'd 914: o_tuple = 10'b1111011010;  // alpha^914
            10'd 915: o_tuple = 10'b1110111101;  // alpha^915
            10'd 916: o_tuple = 10'b1101110011;  // alpha^916
            10'd 917: o_tuple = 10'b1011101111;  // alpha^917
            10'd 918: o_tuple = 10'b0111010111;  // alpha^918
            10'd 919: o_tuple = 10'b1110101110;  // alpha^919
            10'd 920: o_tuple = 10'b1101010101;  // alpha^920
            10'd 921: o_tuple = 10'b1010100011;  // alpha^921
            10'd 922: o_tuple = 10'b0101001111;  // alpha^922
            10'd 923: o_tuple = 10'b1010011110;  // alpha^923
            10'd 924: o_tuple = 10'b0100110101;  // alpha^924
            10'd 925: o_tuple = 10'b1001101010;  // alpha^925
            10'd 926: o_tuple = 10'b0011011101;  // alpha^926
            10'd 927: o_tuple = 10'b0110111010;  // alpha^927
            10'd 928: o_tuple = 10'b1101110100;  // alpha^928
            10'd 929: o_tuple = 10'b1011100001;  // alpha^929
            10'd 930: o_tuple = 10'b0111001011;  // alpha^930
            10'd 931: o_tuple = 10'b1110010110;  // alpha^931
            10'd 932: o_tuple = 10'b1100100101;  // alpha^932
            10'd 933: o_tuple = 10'b1001000011;  // alpha^933
            10'd 934: o_tuple = 10'b0010001111;  // alpha^934
            10'd 935: o_tuple = 10'b0100011110;  // alpha^935
            10'd 936: o_tuple = 10'b1000111100;  // alpha^936
            10'd 937: o_tuple = 10'b0001110001;  // alpha^937
            10'd 938: o_tuple = 10'b0011100010;  // alpha^938
            10'd 939: o_tuple = 10'b0111000100;  // alpha^939
            10'd 940: o_tuple = 10'b1110001000;  // alpha^940
            10'd 941: o_tuple = 10'b1100011001;  // alpha^941
            10'd 942: o_tuple = 10'b1000111011;  // alpha^942
            10'd 943: o_tuple = 10'b0001111111;  // alpha^943
            10'd 944: o_tuple = 10'b0011111110;  // alpha^944
            10'd 945: o_tuple = 10'b0111111100;  // alpha^945
            10'd 946: o_tuple = 10'b1111111000;  // alpha^946
            10'd 947: o_tuple = 10'b1111111001;  // alpha^947
            10'd 948: o_tuple = 10'b1111111011;  // alpha^948
            10'd 949: o_tuple = 10'b1111111111;  // alpha^949
            10'd 950: o_tuple = 10'b1111110111;  // alpha^950
            10'd 951: o_tuple = 10'b1111100111;  // alpha^951
            10'd 952: o_tuple = 10'b1111000111;  // alpha^952
            10'd 953: o_tuple = 10'b1110000111;  // alpha^953
            10'd 954: o_tuple = 10'b1100000111;  // alpha^954
            10'd 955: o_tuple = 10'b1000000111;  // alpha^955
            10'd 956: o_tuple = 10'b0000000111;  // alpha^956
            10'd 957: o_tuple = 10'b0000001110;  // alpha^957
            10'd 958: o_tuple = 10'b0000011100;  // alpha^958
            10'd 959: o_tuple = 10'b0000111000;  // alpha^959
            10'd 960: o_tuple = 10'b0001110000;  // alpha^960
            10'd 961: o_tuple = 10'b0011100000;  // alpha^961
            10'd 962: o_tuple = 10'b0111000000;  // alpha^962
            10'd 963: o_tuple = 10'b1110000000;  // alpha^963
            10'd 964: o_tuple = 10'b1100001001;  // alpha^964
            10'd 965: o_tuple = 10'b1000011011;  // alpha^965
            10'd 966: o_tuple = 10'b0000111111;  // alpha^966
            10'd 967: o_tuple = 10'b0001111110;  // alpha^967
            10'd 968: o_tuple = 10'b0011111100;  // alpha^968
            10'd 969: o_tuple = 10'b0111111000;  // alpha^969
            10'd 970: o_tuple = 10'b1111110000;  // alpha^970
            10'd 971: o_tuple = 10'b1111101001;  // alpha^971
            10'd 972: o_tuple = 10'b1111011011;  // alpha^972
            10'd 973: o_tuple = 10'b1110111111;  // alpha^973
            10'd 974: o_tuple = 10'b1101110111;  // alpha^974
            10'd 975: o_tuple = 10'b1011100111;  // alpha^975
            10'd 976: o_tuple = 10'b0111000111;  // alpha^976
            10'd 977: o_tuple = 10'b1110001110;  // alpha^977
            10'd 978: o_tuple = 10'b1100010101;  // alpha^978
            10'd 979: o_tuple = 10'b1000100011;  // alpha^979
            10'd 980: o_tuple = 10'b0001001111;  // alpha^980
            10'd 981: o_tuple = 10'b0010011110;  // alpha^981
            10'd 982: o_tuple = 10'b0100111100;  // alpha^982
            10'd 983: o_tuple = 10'b1001111000;  // alpha^983
            10'd 984: o_tuple = 10'b0011111001;  // alpha^984
            10'd 985: o_tuple = 10'b0111110010;  // alpha^985
            10'd 986: o_tuple = 10'b1111100100;  // alpha^986
            10'd 987: o_tuple = 10'b1111000001;  // alpha^987
            10'd 988: o_tuple = 10'b1110001011;  // alpha^988
            10'd 989: o_tuple = 10'b1100011111;  // alpha^989
            10'd 990: o_tuple = 10'b1000110111;  // alpha^990
            10'd 991: o_tuple = 10'b0001100111;  // alpha^991
            10'd 992: o_tuple = 10'b0011001110;  // alpha^992
            10'd 993: o_tuple = 10'b0110011100;  // alpha^993
            10'd 994: o_tuple = 10'b1100111000;  // alpha^994
            10'd 995: o_tuple = 10'b1001111001;  // alpha^995
            10'd 996: o_tuple = 10'b0011111011;  // alpha^996
            10'd 997: o_tuple = 10'b0111110110;  // alpha^997
            10'd 998: o_tuple = 10'b1111101100;  // alpha^998
            10'd 999: o_tuple = 10'b1111010001;  // alpha^999
            10'd1000: o_tuple = 10'b1110101011;  // alpha^1000
            10'd1001: o_tuple = 10'b1101011111;  // alpha^1001
            10'd1002: o_tuple = 10'b1010110111;  // alpha^1002
            10'd1003: o_tuple = 10'b0101100111;  // alpha^1003
            10'd1004: o_tuple = 10'b1011001110;  // alpha^1004
            10'd1005: o_tuple = 10'b0110010101;  // alpha^1005
            10'd1006: o_tuple = 10'b1100101010;  // alpha^1006
            10'd1007: o_tuple = 10'b1001011101;  // alpha^1007
            10'd1008: o_tuple = 10'b0010110011;  // alpha^1008
            10'd1009: o_tuple = 10'b0101100110;  // alpha^1009
            10'd1010: o_tuple = 10'b1011001100;  // alpha^1010
            10'd1011: o_tuple = 10'b0110010001;  // alpha^1011
            10'd1012: o_tuple = 10'b1100100010;  // alpha^1012
            10'd1013: o_tuple = 10'b1001001101;  // alpha^1013
            10'd1014: o_tuple = 10'b0010010011;  // alpha^1014
            10'd1015: o_tuple = 10'b0100100110;  // alpha^1015
            10'd1016: o_tuple = 10'b1001001100;  // alpha^1016
            10'd1017: o_tuple = 10'b0010010001;  // alpha^1017
            10'd1018: o_tuple = 10'b0100100010;  // alpha^1018
            10'd1019: o_tuple = 10'b1001000100;  // alpha^1019
            10'd1020: o_tuple = 10'b0010000001;  // alpha^1020
            10'd1021: o_tuple = 10'b0100000010;  // alpha^1021
            10'd1022: o_tuple = 10'b1000000100;  // alpha^1022
            default: o_tuple = 10'd1023;  // Default to zero
        endcase
    end

endmodule


module tuple_to_power_1023_1015(
    input  [9:0] i_tuple,
    output reg [9:0] o_power
);

    always @(*) begin
        case (i_tuple)
            10'b0000000000: o_power = 10'd1023;  // ZERO (power = -1)

            10'b0000000001: o_power = 10'd   0;  // alpha^0
            10'b0000000010: o_power = 10'd   1;  // alpha^1
            10'b0000000100: o_power = 10'd   2;  // alpha^2
            10'b0000001000: o_power = 10'd   3;  // alpha^3
            10'b0000010000: o_power = 10'd   4;  // alpha^4
            10'b0000100000: o_power = 10'd   5;  // alpha^5
            10'b0001000000: o_power = 10'd   6;  // alpha^6
            10'b0010000000: o_power = 10'd   7;  // alpha^7
            10'b0100000000: o_power = 10'd   8;  // alpha^8
            10'b1000000000: o_power = 10'd   9;  // alpha^9
            10'b0000001001: o_power = 10'd  10;  // alpha^10
            10'b0000010010: o_power = 10'd  11;  // alpha^11
            10'b0000100100: o_power = 10'd  12;  // alpha^12
            10'b0001001000: o_power = 10'd  13;  // alpha^13
            10'b0010010000: o_power = 10'd  14;  // alpha^14
            10'b0100100000: o_power = 10'd  15;  // alpha^15
            10'b1001000000: o_power = 10'd  16;  // alpha^16
            10'b0010001001: o_power = 10'd  17;  // alpha^17
            10'b0100010010: o_power = 10'd  18;  // alpha^18
            10'b1000100100: o_power = 10'd  19;  // alpha^19
            10'b0001000001: o_power = 10'd  20;  // alpha^20
            10'b0010000010: o_power = 10'd  21;  // alpha^21
            10'b0100000100: o_power = 10'd  22;  // alpha^22
            10'b1000001000: o_power = 10'd  23;  // alpha^23
            10'b0000011001: o_power = 10'd  24;  // alpha^24
            10'b0000110010: o_power = 10'd  25;  // alpha^25
            10'b0001100100: o_power = 10'd  26;  // alpha^26
            10'b0011001000: o_power = 10'd  27;  // alpha^27
            10'b0110010000: o_power = 10'd  28;  // alpha^28
            10'b1100100000: o_power = 10'd  29;  // alpha^29
            10'b1001001001: o_power = 10'd  30;  // alpha^30
            10'b0010011011: o_power = 10'd  31;  // alpha^31
            10'b0100110110: o_power = 10'd  32;  // alpha^32
            10'b1001101100: o_power = 10'd  33;  // alpha^33
            10'b0011010001: o_power = 10'd  34;  // alpha^34
            10'b0110100010: o_power = 10'd  35;  // alpha^35
            10'b1101000100: o_power = 10'd  36;  // alpha^36
            10'b1010000001: o_power = 10'd  37;  // alpha^37
            10'b0100001011: o_power = 10'd  38;  // alpha^38
            10'b1000010110: o_power = 10'd  39;  // alpha^39
            10'b0000100101: o_power = 10'd  40;  // alpha^40
            10'b0001001010: o_power = 10'd  41;  // alpha^41
            10'b0010010100: o_power = 10'd  42;  // alpha^42
            10'b0100101000: o_power = 10'd  43;  // alpha^43
            10'b1001010000: o_power = 10'd  44;  // alpha^44
            10'b0010101001: o_power = 10'd  45;  // alpha^45
            10'b0101010010: o_power = 10'd  46;  // alpha^46
            10'b1010100100: o_power = 10'd  47;  // alpha^47
            10'b0101000001: o_power = 10'd  48;  // alpha^48
            10'b1010000010: o_power = 10'd  49;  // alpha^49
            10'b0100001101: o_power = 10'd  50;  // alpha^50
            10'b1000011010: o_power = 10'd  51;  // alpha^51
            10'b0000111101: o_power = 10'd  52;  // alpha^52
            10'b0001111010: o_power = 10'd  53;  // alpha^53
            10'b0011110100: o_power = 10'd  54;  // alpha^54
            10'b0111101000: o_power = 10'd  55;  // alpha^55
            10'b1111010000: o_power = 10'd  56;  // alpha^56
            10'b1110101001: o_power = 10'd  57;  // alpha^57
            10'b1101011011: o_power = 10'd  58;  // alpha^58
            10'b1010111111: o_power = 10'd  59;  // alpha^59
            10'b0101110111: o_power = 10'd  60;  // alpha^60
            10'b1011101110: o_power = 10'd  61;  // alpha^61
            10'b0111010101: o_power = 10'd  62;  // alpha^62
            10'b1110101010: o_power = 10'd  63;  // alpha^63
            10'b1101011101: o_power = 10'd  64;  // alpha^64
            10'b1010110011: o_power = 10'd  65;  // alpha^65
            10'b0101101111: o_power = 10'd  66;  // alpha^66
            10'b1011011110: o_power = 10'd  67;  // alpha^67
            10'b0110110101: o_power = 10'd  68;  // alpha^68
            10'b1101101010: o_power = 10'd  69;  // alpha^69
            10'b1011011101: o_power = 10'd  70;  // alpha^70
            10'b0110110011: o_power = 10'd  71;  // alpha^71
            10'b1101100110: o_power = 10'd  72;  // alpha^72
            10'b1011000101: o_power = 10'd  73;  // alpha^73
            10'b0110000011: o_power = 10'd  74;  // alpha^74
            10'b1100000110: o_power = 10'd  75;  // alpha^75
            10'b1000000101: o_power = 10'd  76;  // alpha^76
            10'b0000000011: o_power = 10'd  77;  // alpha^77
            10'b0000000110: o_power = 10'd  78;  // alpha^78
            10'b0000001100: o_power = 10'd  79;  // alpha^79
            10'b0000011000: o_power = 10'd  80;  // alpha^80
            10'b0000110000: o_power = 10'd  81;  // alpha^81
            10'b0001100000: o_power = 10'd  82;  // alpha^82
            10'b0011000000: o_power = 10'd  83;  // alpha^83
            10'b0110000000: o_power = 10'd  84;  // alpha^84
            10'b1100000000: o_power = 10'd  85;  // alpha^85
            10'b1000001001: o_power = 10'd  86;  // alpha^86
            10'b0000011011: o_power = 10'd  87;  // alpha^87
            10'b0000110110: o_power = 10'd  88;  // alpha^88
            10'b0001101100: o_power = 10'd  89;  // alpha^89
            10'b0011011000: o_power = 10'd  90;  // alpha^90
            10'b0110110000: o_power = 10'd  91;  // alpha^91
            10'b1101100000: o_power = 10'd  92;  // alpha^92
            10'b1011001001: o_power = 10'd  93;  // alpha^93
            10'b0110011011: o_power = 10'd  94;  // alpha^94
            10'b1100110110: o_power = 10'd  95;  // alpha^95
            10'b1001100101: o_power = 10'd  96;  // alpha^96
            10'b0011000011: o_power = 10'd  97;  // alpha^97
            10'b0110000110: o_power = 10'd  98;  // alpha^98
            10'b1100001100: o_power = 10'd  99;  // alpha^99
            10'b1000010001: o_power = 10'd 100;  // alpha^100
            10'b0000101011: o_power = 10'd 101;  // alpha^101
            10'b0001010110: o_power = 10'd 102;  // alpha^102
            10'b0010101100: o_power = 10'd 103;  // alpha^103
            10'b0101011000: o_power = 10'd 104;  // alpha^104
            10'b1010110000: o_power = 10'd 105;  // alpha^105
            10'b0101101001: o_power = 10'd 106;  // alpha^106
            10'b1011010010: o_power = 10'd 107;  // alpha^107
            10'b0110101101: o_power = 10'd 108;  // alpha^108
            10'b1101011010: o_power = 10'd 109;  // alpha^109
            10'b1010111101: o_power = 10'd 110;  // alpha^110
            10'b0101110011: o_power = 10'd 111;  // alpha^111
            10'b1011100110: o_power = 10'd 112;  // alpha^112
            10'b0111000101: o_power = 10'd 113;  // alpha^113
            10'b1110001010: o_power = 10'd 114;  // alpha^114
            10'b1100011101: o_power = 10'd 115;  // alpha^115
            10'b1000110011: o_power = 10'd 116;  // alpha^116
            10'b0001101111: o_power = 10'd 117;  // alpha^117
            10'b0011011110: o_power = 10'd 118;  // alpha^118
            10'b0110111100: o_power = 10'd 119;  // alpha^119
            10'b1101111000: o_power = 10'd 120;  // alpha^120
            10'b1011111001: o_power = 10'd 121;  // alpha^121
            10'b0111111011: o_power = 10'd 122;  // alpha^122
            10'b1111110110: o_power = 10'd 123;  // alpha^123
            10'b1111100101: o_power = 10'd 124;  // alpha^124
            10'b1111000011: o_power = 10'd 125;  // alpha^125
            10'b1110001111: o_power = 10'd 126;  // alpha^126
            10'b1100010111: o_power = 10'd 127;  // alpha^127
            10'b1000100111: o_power = 10'd 128;  // alpha^128
            10'b0001000111: o_power = 10'd 129;  // alpha^129
            10'b0010001110: o_power = 10'd 130;  // alpha^130
            10'b0100011100: o_power = 10'd 131;  // alpha^131
            10'b1000111000: o_power = 10'd 132;  // alpha^132
            10'b0001111001: o_power = 10'd 133;  // alpha^133
            10'b0011110010: o_power = 10'd 134;  // alpha^134
            10'b0111100100: o_power = 10'd 135;  // alpha^135
            10'b1111001000: o_power = 10'd 136;  // alpha^136
            10'b1110011001: o_power = 10'd 137;  // alpha^137
            10'b1100111011: o_power = 10'd 138;  // alpha^138
            10'b1001111111: o_power = 10'd 139;  // alpha^139
            10'b0011110111: o_power = 10'd 140;  // alpha^140
            10'b0111101110: o_power = 10'd 141;  // alpha^141
            10'b1111011100: o_power = 10'd 142;  // alpha^142
            10'b1110110001: o_power = 10'd 143;  // alpha^143
            10'b1101101011: o_power = 10'd 144;  // alpha^144
            10'b1011011111: o_power = 10'd 145;  // alpha^145
            10'b0110110111: o_power = 10'd 146;  // alpha^146
            10'b1101101110: o_power = 10'd 147;  // alpha^147
            10'b1011010101: o_power = 10'd 148;  // alpha^148
            10'b0110100011: o_power = 10'd 149;  // alpha^149
            10'b1101000110: o_power = 10'd 150;  // alpha^150
            10'b1010000101: o_power = 10'd 151;  // alpha^151
            10'b0100000011: o_power = 10'd 152;  // alpha^152
            10'b1000000110: o_power = 10'd 153;  // alpha^153
            10'b0000000101: o_power = 10'd 154;  // alpha^154
            10'b0000001010: o_power = 10'd 155;  // alpha^155
            10'b0000010100: o_power = 10'd 156;  // alpha^156
            10'b0000101000: o_power = 10'd 157;  // alpha^157
            10'b0001010000: o_power = 10'd 158;  // alpha^158
            10'b0010100000: o_power = 10'd 159;  // alpha^159
            10'b0101000000: o_power = 10'd 160;  // alpha^160
            10'b1010000000: o_power = 10'd 161;  // alpha^161
            10'b0100001001: o_power = 10'd 162;  // alpha^162
            10'b1000010010: o_power = 10'd 163;  // alpha^163
            10'b0000101101: o_power = 10'd 164;  // alpha^164
            10'b0001011010: o_power = 10'd 165;  // alpha^165
            10'b0010110100: o_power = 10'd 166;  // alpha^166
            10'b0101101000: o_power = 10'd 167;  // alpha^167
            10'b1011010000: o_power = 10'd 168;  // alpha^168
            10'b0110101001: o_power = 10'd 169;  // alpha^169
            10'b1101010010: o_power = 10'd 170;  // alpha^170
            10'b1010101101: o_power = 10'd 171;  // alpha^171
            10'b0101010011: o_power = 10'd 172;  // alpha^172
            10'b1010100110: o_power = 10'd 173;  // alpha^173
            10'b0101000101: o_power = 10'd 174;  // alpha^174
            10'b1010001010: o_power = 10'd 175;  // alpha^175
            10'b0100011101: o_power = 10'd 176;  // alpha^176
            10'b1000111010: o_power = 10'd 177;  // alpha^177
            10'b0001111101: o_power = 10'd 178;  // alpha^178
            10'b0011111010: o_power = 10'd 179;  // alpha^179
            10'b0111110100: o_power = 10'd 180;  // alpha^180
            10'b1111101000: o_power = 10'd 181;  // alpha^181
            10'b1111011001: o_power = 10'd 182;  // alpha^182
            10'b1110111011: o_power = 10'd 183;  // alpha^183
            10'b1101111111: o_power = 10'd 184;  // alpha^184
            10'b1011110111: o_power = 10'd 185;  // alpha^185
            10'b0111100111: o_power = 10'd 186;  // alpha^186
            10'b1111001110: o_power = 10'd 187;  // alpha^187
            10'b1110010101: o_power = 10'd 188;  // alpha^188
            10'b1100100011: o_power = 10'd 189;  // alpha^189
            10'b1001001111: o_power = 10'd 190;  // alpha^190
            10'b0010010111: o_power = 10'd 191;  // alpha^191
            10'b0100101110: o_power = 10'd 192;  // alpha^192
            10'b1001011100: o_power = 10'd 193;  // alpha^193
            10'b0010110001: o_power = 10'd 194;  // alpha^194
            10'b0101100010: o_power = 10'd 195;  // alpha^195
            10'b1011000100: o_power = 10'd 196;  // alpha^196
            10'b0110000001: o_power = 10'd 197;  // alpha^197
            10'b1100000010: o_power = 10'd 198;  // alpha^198
            10'b1000001101: o_power = 10'd 199;  // alpha^199
            10'b0000010011: o_power = 10'd 200;  // alpha^200
            10'b0000100110: o_power = 10'd 201;  // alpha^201
            10'b0001001100: o_power = 10'd 202;  // alpha^202
            10'b0010011000: o_power = 10'd 203;  // alpha^203
            10'b0100110000: o_power = 10'd 204;  // alpha^204
            10'b1001100000: o_power = 10'd 205;  // alpha^205
            10'b0011001001: o_power = 10'd 206;  // alpha^206
            10'b0110010010: o_power = 10'd 207;  // alpha^207
            10'b1100100100: o_power = 10'd 208;  // alpha^208
            10'b1001000001: o_power = 10'd 209;  // alpha^209
            10'b0010001011: o_power = 10'd 210;  // alpha^210
            10'b0100010110: o_power = 10'd 211;  // alpha^211
            10'b1000101100: o_power = 10'd 212;  // alpha^212
            10'b0001010001: o_power = 10'd 213;  // alpha^213
            10'b0010100010: o_power = 10'd 214;  // alpha^214
            10'b0101000100: o_power = 10'd 215;  // alpha^215
            10'b1010001000: o_power = 10'd 216;  // alpha^216
            10'b0100011001: o_power = 10'd 217;  // alpha^217
            10'b1000110010: o_power = 10'd 218;  // alpha^218
            10'b0001101101: o_power = 10'd 219;  // alpha^219
            10'b0011011010: o_power = 10'd 220;  // alpha^220
            10'b0110110100: o_power = 10'd 221;  // alpha^221
            10'b1101101000: o_power = 10'd 222;  // alpha^222
            10'b1011011001: o_power = 10'd 223;  // alpha^223
            10'b0110111011: o_power = 10'd 224;  // alpha^224
            10'b1101110110: o_power = 10'd 225;  // alpha^225
            10'b1011100101: o_power = 10'd 226;  // alpha^226
            10'b0111000011: o_power = 10'd 227;  // alpha^227
            10'b1110000110: o_power = 10'd 228;  // alpha^228
            10'b1100000101: o_power = 10'd 229;  // alpha^229
            10'b1000000011: o_power = 10'd 230;  // alpha^230
            10'b0000001111: o_power = 10'd 231;  // alpha^231
            10'b0000011110: o_power = 10'd 232;  // alpha^232
            10'b0000111100: o_power = 10'd 233;  // alpha^233
            10'b0001111000: o_power = 10'd 234;  // alpha^234
            10'b0011110000: o_power = 10'd 235;  // alpha^235
            10'b0111100000: o_power = 10'd 236;  // alpha^236
            10'b1111000000: o_power = 10'd 237;  // alpha^237
            10'b1110001001: o_power = 10'd 238;  // alpha^238
            10'b1100011011: o_power = 10'd 239;  // alpha^239
            10'b1000111111: o_power = 10'd 240;  // alpha^240
            10'b0001110111: o_power = 10'd 241;  // alpha^241
            10'b0011101110: o_power = 10'd 242;  // alpha^242
            10'b0111011100: o_power = 10'd 243;  // alpha^243
            10'b1110111000: o_power = 10'd 244;  // alpha^244
            10'b1101111001: o_power = 10'd 245;  // alpha^245
            10'b1011111011: o_power = 10'd 246;  // alpha^246
            10'b0111111111: o_power = 10'd 247;  // alpha^247
            10'b1111111110: o_power = 10'd 248;  // alpha^248
            10'b1111110101: o_power = 10'd 249;  // alpha^249
            10'b1111100011: o_power = 10'd 250;  // alpha^250
            10'b1111001111: o_power = 10'd 251;  // alpha^251
            10'b1110010111: o_power = 10'd 252;  // alpha^252
            10'b1100100111: o_power = 10'd 253;  // alpha^253
            10'b1001000111: o_power = 10'd 254;  // alpha^254
            10'b0010000111: o_power = 10'd 255;  // alpha^255
            10'b0100001110: o_power = 10'd 256;  // alpha^256
            10'b1000011100: o_power = 10'd 257;  // alpha^257
            10'b0000110001: o_power = 10'd 258;  // alpha^258
            10'b0001100010: o_power = 10'd 259;  // alpha^259
            10'b0011000100: o_power = 10'd 260;  // alpha^260
            10'b0110001000: o_power = 10'd 261;  // alpha^261
            10'b1100010000: o_power = 10'd 262;  // alpha^262
            10'b1000101001: o_power = 10'd 263;  // alpha^263
            10'b0001011011: o_power = 10'd 264;  // alpha^264
            10'b0010110110: o_power = 10'd 265;  // alpha^265
            10'b0101101100: o_power = 10'd 266;  // alpha^266
            10'b1011011000: o_power = 10'd 267;  // alpha^267
            10'b0110111001: o_power = 10'd 268;  // alpha^268
            10'b1101110010: o_power = 10'd 269;  // alpha^269
            10'b1011101101: o_power = 10'd 270;  // alpha^270
            10'b0111010011: o_power = 10'd 271;  // alpha^271
            10'b1110100110: o_power = 10'd 272;  // alpha^272
            10'b1101000101: o_power = 10'd 273;  // alpha^273
            10'b1010000011: o_power = 10'd 274;  // alpha^274
            10'b0100001111: o_power = 10'd 275;  // alpha^275
            10'b1000011110: o_power = 10'd 276;  // alpha^276
            10'b0000110101: o_power = 10'd 277;  // alpha^277
            10'b0001101010: o_power = 10'd 278;  // alpha^278
            10'b0011010100: o_power = 10'd 279;  // alpha^279
            10'b0110101000: o_power = 10'd 280;  // alpha^280
            10'b1101010000: o_power = 10'd 281;  // alpha^281
            10'b1010101001: o_power = 10'd 282;  // alpha^282
            10'b0101011011: o_power = 10'd 283;  // alpha^283
            10'b1010110110: o_power = 10'd 284;  // alpha^284
            10'b0101100101: o_power = 10'd 285;  // alpha^285
            10'b1011001010: o_power = 10'd 286;  // alpha^286
            10'b0110011101: o_power = 10'd 287;  // alpha^287
            10'b1100111010: o_power = 10'd 288;  // alpha^288
            10'b1001111101: o_power = 10'd 289;  // alpha^289
            10'b0011110011: o_power = 10'd 290;  // alpha^290
            10'b0111100110: o_power = 10'd 291;  // alpha^291
            10'b1111001100: o_power = 10'd 292;  // alpha^292
            10'b1110010001: o_power = 10'd 293;  // alpha^293
            10'b1100101011: o_power = 10'd 294;  // alpha^294
            10'b1001011111: o_power = 10'd 295;  // alpha^295
            10'b0010110111: o_power = 10'd 296;  // alpha^296
            10'b0101101110: o_power = 10'd 297;  // alpha^297
            10'b1011011100: o_power = 10'd 298;  // alpha^298
            10'b0110110001: o_power = 10'd 299;  // alpha^299
            10'b1101100010: o_power = 10'd 300;  // alpha^300
            10'b1011001101: o_power = 10'd 301;  // alpha^301
            10'b0110010011: o_power = 10'd 302;  // alpha^302
            10'b1100100110: o_power = 10'd 303;  // alpha^303
            10'b1001000101: o_power = 10'd 304;  // alpha^304
            10'b0010000011: o_power = 10'd 305;  // alpha^305
            10'b0100000110: o_power = 10'd 306;  // alpha^306
            10'b1000001100: o_power = 10'd 307;  // alpha^307
            10'b0000010001: o_power = 10'd 308;  // alpha^308
            10'b0000100010: o_power = 10'd 309;  // alpha^309
            10'b0001000100: o_power = 10'd 310;  // alpha^310
            10'b0010001000: o_power = 10'd 311;  // alpha^311
            10'b0100010000: o_power = 10'd 312;  // alpha^312
            10'b1000100000: o_power = 10'd 313;  // alpha^313
            10'b0001001001: o_power = 10'd 314;  // alpha^314
            10'b0010010010: o_power = 10'd 315;  // alpha^315
            10'b0100100100: o_power = 10'd 316;  // alpha^316
            10'b1001001000: o_power = 10'd 317;  // alpha^317
            10'b0010011001: o_power = 10'd 318;  // alpha^318
            10'b0100110010: o_power = 10'd 319;  // alpha^319
            10'b1001100100: o_power = 10'd 320;  // alpha^320
            10'b0011000001: o_power = 10'd 321;  // alpha^321
            10'b0110000010: o_power = 10'd 322;  // alpha^322
            10'b1100000100: o_power = 10'd 323;  // alpha^323
            10'b1000000001: o_power = 10'd 324;  // alpha^324
            10'b0000001011: o_power = 10'd 325;  // alpha^325
            10'b0000010110: o_power = 10'd 326;  // alpha^326
            10'b0000101100: o_power = 10'd 327;  // alpha^327
            10'b0001011000: o_power = 10'd 328;  // alpha^328
            10'b0010110000: o_power = 10'd 329;  // alpha^329
            10'b0101100000: o_power = 10'd 330;  // alpha^330
            10'b1011000000: o_power = 10'd 331;  // alpha^331
            10'b0110001001: o_power = 10'd 332;  // alpha^332
            10'b1100010010: o_power = 10'd 333;  // alpha^333
            10'b1000101101: o_power = 10'd 334;  // alpha^334
            10'b0001010011: o_power = 10'd 335;  // alpha^335
            10'b0010100110: o_power = 10'd 336;  // alpha^336
            10'b0101001100: o_power = 10'd 337;  // alpha^337
            10'b1010011000: o_power = 10'd 338;  // alpha^338
            10'b0100111001: o_power = 10'd 339;  // alpha^339
            10'b1001110010: o_power = 10'd 340;  // alpha^340
            10'b0011101101: o_power = 10'd 341;  // alpha^341
            10'b0111011010: o_power = 10'd 342;  // alpha^342
            10'b1110110100: o_power = 10'd 343;  // alpha^343
            10'b1101100001: o_power = 10'd 344;  // alpha^344
            10'b1011001011: o_power = 10'd 345;  // alpha^345
            10'b0110011111: o_power = 10'd 346;  // alpha^346
            10'b1100111110: o_power = 10'd 347;  // alpha^347
            10'b1001110101: o_power = 10'd 348;  // alpha^348
            10'b0011100011: o_power = 10'd 349;  // alpha^349
            10'b0111000110: o_power = 10'd 350;  // alpha^350
            10'b1110001100: o_power = 10'd 351;  // alpha^351
            10'b1100010001: o_power = 10'd 352;  // alpha^352
            10'b1000101011: o_power = 10'd 353;  // alpha^353
            10'b0001011111: o_power = 10'd 354;  // alpha^354
            10'b0010111110: o_power = 10'd 355;  // alpha^355
            10'b0101111100: o_power = 10'd 356;  // alpha^356
            10'b1011111000: o_power = 10'd 357;  // alpha^357
            10'b0111111001: o_power = 10'd 358;  // alpha^358
            10'b1111110010: o_power = 10'd 359;  // alpha^359
            10'b1111101101: o_power = 10'd 360;  // alpha^360
            10'b1111010011: o_power = 10'd 361;  // alpha^361
            10'b1110101111: o_power = 10'd 362;  // alpha^362
            10'b1101010111: o_power = 10'd 363;  // alpha^363
            10'b1010100111: o_power = 10'd 364;  // alpha^364
            10'b0101000111: o_power = 10'd 365;  // alpha^365
            10'b1010001110: o_power = 10'd 366;  // alpha^366
            10'b0100010101: o_power = 10'd 367;  // alpha^367
            10'b1000101010: o_power = 10'd 368;  // alpha^368
            10'b0001011101: o_power = 10'd 369;  // alpha^369
            10'b0010111010: o_power = 10'd 370;  // alpha^370
            10'b0101110100: o_power = 10'd 371;  // alpha^371
            10'b1011101000: o_power = 10'd 372;  // alpha^372
            10'b0111011001: o_power = 10'd 373;  // alpha^373
            10'b1110110010: o_power = 10'd 374;  // alpha^374
            10'b1101101101: o_power = 10'd 375;  // alpha^375
            10'b1011010011: o_power = 10'd 376;  // alpha^376
            10'b0110101111: o_power = 10'd 377;  // alpha^377
            10'b1101011110: o_power = 10'd 378;  // alpha^378
            10'b1010110101: o_power = 10'd 379;  // alpha^379
            10'b0101100011: o_power = 10'd 380;  // alpha^380
            10'b1011000110: o_power = 10'd 381;  // alpha^381
            10'b0110000101: o_power = 10'd 382;  // alpha^382
            10'b1100001010: o_power = 10'd 383;  // alpha^383
            10'b1000011101: o_power = 10'd 384;  // alpha^384
            10'b0000110011: o_power = 10'd 385;  // alpha^385
            10'b0001100110: o_power = 10'd 386;  // alpha^386
            10'b0011001100: o_power = 10'd 387;  // alpha^387
            10'b0110011000: o_power = 10'd 388;  // alpha^388
            10'b1100110000: o_power = 10'd 389;  // alpha^389
            10'b1001101001: o_power = 10'd 390;  // alpha^390
            10'b0011011011: o_power = 10'd 391;  // alpha^391
            10'b0110110110: o_power = 10'd 392;  // alpha^392
            10'b1101101100: o_power = 10'd 393;  // alpha^393
            10'b1011010001: o_power = 10'd 394;  // alpha^394
            10'b0110101011: o_power = 10'd 395;  // alpha^395
            10'b1101010110: o_power = 10'd 396;  // alpha^396
            10'b1010100101: o_power = 10'd 397;  // alpha^397
            10'b0101000011: o_power = 10'd 398;  // alpha^398
            10'b1010000110: o_power = 10'd 399;  // alpha^399
            10'b0100000101: o_power = 10'd 400;  // alpha^400
            10'b1000001010: o_power = 10'd 401;  // alpha^401
            10'b0000011101: o_power = 10'd 402;  // alpha^402
            10'b0000111010: o_power = 10'd 403;  // alpha^403
            10'b0001110100: o_power = 10'd 404;  // alpha^404
            10'b0011101000: o_power = 10'd 405;  // alpha^405
            10'b0111010000: o_power = 10'd 406;  // alpha^406
            10'b1110100000: o_power = 10'd 407;  // alpha^407
            10'b1101001001: o_power = 10'd 408;  // alpha^408
            10'b1010011011: o_power = 10'd 409;  // alpha^409
            10'b0100111111: o_power = 10'd 410;  // alpha^410
            10'b1001111110: o_power = 10'd 411;  // alpha^411
            10'b0011110101: o_power = 10'd 412;  // alpha^412
            10'b0111101010: o_power = 10'd 413;  // alpha^413
            10'b1111010100: o_power = 10'd 414;  // alpha^414
            10'b1110100001: o_power = 10'd 415;  // alpha^415
            10'b1101001011: o_power = 10'd 416;  // alpha^416
            10'b1010011111: o_power = 10'd 417;  // alpha^417
            10'b0100110111: o_power = 10'd 418;  // alpha^418
            10'b1001101110: o_power = 10'd 419;  // alpha^419
            10'b0011010101: o_power = 10'd 420;  // alpha^420
            10'b0110101010: o_power = 10'd 421;  // alpha^421
            10'b1101010100: o_power = 10'd 422;  // alpha^422
            10'b1010100001: o_power = 10'd 423;  // alpha^423
            10'b0101001011: o_power = 10'd 424;  // alpha^424
            10'b1010010110: o_power = 10'd 425;  // alpha^425
            10'b0100100101: o_power = 10'd 426;  // alpha^426
            10'b1001001010: o_power = 10'd 427;  // alpha^427
            10'b0010011101: o_power = 10'd 428;  // alpha^428
            10'b0100111010: o_power = 10'd 429;  // alpha^429
            10'b1001110100: o_power = 10'd 430;  // alpha^430
            10'b0011100001: o_power = 10'd 431;  // alpha^431
            10'b0111000010: o_power = 10'd 432;  // alpha^432
            10'b1110000100: o_power = 10'd 433;  // alpha^433
            10'b1100000001: o_power = 10'd 434;  // alpha^434
            10'b1000001011: o_power = 10'd 435;  // alpha^435
            10'b0000011111: o_power = 10'd 436;  // alpha^436
            10'b0000111110: o_power = 10'd 437;  // alpha^437
            10'b0001111100: o_power = 10'd 438;  // alpha^438
            10'b0011111000: o_power = 10'd 439;  // alpha^439
            10'b0111110000: o_power = 10'd 440;  // alpha^440
            10'b1111100000: o_power = 10'd 441;  // alpha^441
            10'b1111001001: o_power = 10'd 442;  // alpha^442
            10'b1110011011: o_power = 10'd 443;  // alpha^443
            10'b1100111111: o_power = 10'd 444;  // alpha^444
            10'b1001110111: o_power = 10'd 445;  // alpha^445
            10'b0011100111: o_power = 10'd 446;  // alpha^446
            10'b0111001110: o_power = 10'd 447;  // alpha^447
            10'b1110011100: o_power = 10'd 448;  // alpha^448
            10'b1100110001: o_power = 10'd 449;  // alpha^449
            10'b1001101011: o_power = 10'd 450;  // alpha^450
            10'b0011011111: o_power = 10'd 451;  // alpha^451
            10'b0110111110: o_power = 10'd 452;  // alpha^452
            10'b1101111100: o_power = 10'd 453;  // alpha^453
            10'b1011110001: o_power = 10'd 454;  // alpha^454
            10'b0111101011: o_power = 10'd 455;  // alpha^455
            10'b1111010110: o_power = 10'd 456;  // alpha^456
            10'b1110100101: o_power = 10'd 457;  // alpha^457
            10'b1101000011: o_power = 10'd 458;  // alpha^458
            10'b1010001111: o_power = 10'd 459;  // alpha^459
            10'b0100010111: o_power = 10'd 460;  // alpha^460
            10'b1000101110: o_power = 10'd 461;  // alpha^461
            10'b0001010101: o_power = 10'd 462;  // alpha^462
            10'b0010101010: o_power = 10'd 463;  // alpha^463
            10'b0101010100: o_power = 10'd 464;  // alpha^464
            10'b1010101000: o_power = 10'd 465;  // alpha^465
            10'b0101011001: o_power = 10'd 466;  // alpha^466
            10'b1010110010: o_power = 10'd 467;  // alpha^467
            10'b0101101101: o_power = 10'd 468;  // alpha^468
            10'b1011011010: o_power = 10'd 469;  // alpha^469
            10'b0110111101: o_power = 10'd 470;  // alpha^470
            10'b1101111010: o_power = 10'd 471;  // alpha^471
            10'b1011111101: o_power = 10'd 472;  // alpha^472
            10'b0111110011: o_power = 10'd 473;  // alpha^473
            10'b1111100110: o_power = 10'd 474;  // alpha^474
            10'b1111000101: o_power = 10'd 475;  // alpha^475
            10'b1110000011: o_power = 10'd 476;  // alpha^476
            10'b1100001111: o_power = 10'd 477;  // alpha^477
            10'b1000010111: o_power = 10'd 478;  // alpha^478
            10'b0000100111: o_power = 10'd 479;  // alpha^479
            10'b0001001110: o_power = 10'd 480;  // alpha^480
            10'b0010011100: o_power = 10'd 481;  // alpha^481
            10'b0100111000: o_power = 10'd 482;  // alpha^482
            10'b1001110000: o_power = 10'd 483;  // alpha^483
            10'b0011101001: o_power = 10'd 484;  // alpha^484
            10'b0111010010: o_power = 10'd 485;  // alpha^485
            10'b1110100100: o_power = 10'd 486;  // alpha^486
            10'b1101000001: o_power = 10'd 487;  // alpha^487
            10'b1010001011: o_power = 10'd 488;  // alpha^488
            10'b0100011111: o_power = 10'd 489;  // alpha^489
            10'b1000111110: o_power = 10'd 490;  // alpha^490
            10'b0001110101: o_power = 10'd 491;  // alpha^491
            10'b0011101010: o_power = 10'd 492;  // alpha^492
            10'b0111010100: o_power = 10'd 493;  // alpha^493
            10'b1110101000: o_power = 10'd 494;  // alpha^494
            10'b1101011001: o_power = 10'd 495;  // alpha^495
            10'b1010111011: o_power = 10'd 496;  // alpha^496
            10'b0101111111: o_power = 10'd 497;  // alpha^497
            10'b1011111110: o_power = 10'd 498;  // alpha^498
            10'b0111110101: o_power = 10'd 499;  // alpha^499
            10'b1111101010: o_power = 10'd 500;  // alpha^500
            10'b1111011101: o_power = 10'd 501;  // alpha^501
            10'b1110110011: o_power = 10'd 502;  // alpha^502
            10'b1101101111: o_power = 10'd 503;  // alpha^503
            10'b1011010111: o_power = 10'd 504;  // alpha^504
            10'b0110100111: o_power = 10'd 505;  // alpha^505
            10'b1101001110: o_power = 10'd 506;  // alpha^506
            10'b1010010101: o_power = 10'd 507;  // alpha^507
            10'b0100100011: o_power = 10'd 508;  // alpha^508
            10'b1001000110: o_power = 10'd 509;  // alpha^509
            10'b0010000101: o_power = 10'd 510;  // alpha^510
            10'b0100001010: o_power = 10'd 511;  // alpha^511
            10'b1000010100: o_power = 10'd 512;  // alpha^512
            10'b0000100001: o_power = 10'd 513;  // alpha^513
            10'b0001000010: o_power = 10'd 514;  // alpha^514
            10'b0010000100: o_power = 10'd 515;  // alpha^515
            10'b0100001000: o_power = 10'd 516;  // alpha^516
            10'b1000010000: o_power = 10'd 517;  // alpha^517
            10'b0000101001: o_power = 10'd 518;  // alpha^518
            10'b0001010010: o_power = 10'd 519;  // alpha^519
            10'b0010100100: o_power = 10'd 520;  // alpha^520
            10'b0101001000: o_power = 10'd 521;  // alpha^521
            10'b1010010000: o_power = 10'd 522;  // alpha^522
            10'b0100101001: o_power = 10'd 523;  // alpha^523
            10'b1001010010: o_power = 10'd 524;  // alpha^524
            10'b0010101101: o_power = 10'd 525;  // alpha^525
            10'b0101011010: o_power = 10'd 526;  // alpha^526
            10'b1010110100: o_power = 10'd 527;  // alpha^527
            10'b0101100001: o_power = 10'd 528;  // alpha^528
            10'b1011000010: o_power = 10'd 529;  // alpha^529
            10'b0110001101: o_power = 10'd 530;  // alpha^530
            10'b1100011010: o_power = 10'd 531;  // alpha^531
            10'b1000111101: o_power = 10'd 532;  // alpha^532
            10'b0001110011: o_power = 10'd 533;  // alpha^533
            10'b0011100110: o_power = 10'd 534;  // alpha^534
            10'b0111001100: o_power = 10'd 535;  // alpha^535
            10'b1110011000: o_power = 10'd 536;  // alpha^536
            10'b1100111001: o_power = 10'd 537;  // alpha^537
            10'b1001111011: o_power = 10'd 538;  // alpha^538
            10'b0011111111: o_power = 10'd 539;  // alpha^539
            10'b0111111110: o_power = 10'd 540;  // alpha^540
            10'b1111111100: o_power = 10'd 541;  // alpha^541
            10'b1111110001: o_power = 10'd 542;  // alpha^542
            10'b1111101011: o_power = 10'd 543;  // alpha^543
            10'b1111011111: o_power = 10'd 544;  // alpha^544
            10'b1110110111: o_power = 10'd 545;  // alpha^545
            10'b1101100111: o_power = 10'd 546;  // alpha^546
            10'b1011000111: o_power = 10'd 547;  // alpha^547
            10'b0110000111: o_power = 10'd 548;  // alpha^548
            10'b1100001110: o_power = 10'd 549;  // alpha^549
            10'b1000010101: o_power = 10'd 550;  // alpha^550
            10'b0000100011: o_power = 10'd 551;  // alpha^551
            10'b0001000110: o_power = 10'd 552;  // alpha^552
            10'b0010001100: o_power = 10'd 553;  // alpha^553
            10'b0100011000: o_power = 10'd 554;  // alpha^554
            10'b1000110000: o_power = 10'd 555;  // alpha^555
            10'b0001101001: o_power = 10'd 556;  // alpha^556
            10'b0011010010: o_power = 10'd 557;  // alpha^557
            10'b0110100100: o_power = 10'd 558;  // alpha^558
            10'b1101001000: o_power = 10'd 559;  // alpha^559
            10'b1010011001: o_power = 10'd 560;  // alpha^560
            10'b0100111011: o_power = 10'd 561;  // alpha^561
            10'b1001110110: o_power = 10'd 562;  // alpha^562
            10'b0011100101: o_power = 10'd 563;  // alpha^563
            10'b0111001010: o_power = 10'd 564;  // alpha^564
            10'b1110010100: o_power = 10'd 565;  // alpha^565
            10'b1100100001: o_power = 10'd 566;  // alpha^566
            10'b1001001011: o_power = 10'd 567;  // alpha^567
            10'b0010011111: o_power = 10'd 568;  // alpha^568
            10'b0100111110: o_power = 10'd 569;  // alpha^569
            10'b1001111100: o_power = 10'd 570;  // alpha^570
            10'b0011110001: o_power = 10'd 571;  // alpha^571
            10'b0111100010: o_power = 10'd 572;  // alpha^572
            10'b1111000100: o_power = 10'd 573;  // alpha^573
            10'b1110000001: o_power = 10'd 574;  // alpha^574
            10'b1100001011: o_power = 10'd 575;  // alpha^575
            10'b1000011111: o_power = 10'd 576;  // alpha^576
            10'b0000110111: o_power = 10'd 577;  // alpha^577
            10'b0001101110: o_power = 10'd 578;  // alpha^578
            10'b0011011100: o_power = 10'd 579;  // alpha^579
            10'b0110111000: o_power = 10'd 580;  // alpha^580
            10'b1101110000: o_power = 10'd 581;  // alpha^581
            10'b1011101001: o_power = 10'd 582;  // alpha^582
            10'b0111011011: o_power = 10'd 583;  // alpha^583
            10'b1110110110: o_power = 10'd 584;  // alpha^584
            10'b1101100101: o_power = 10'd 585;  // alpha^585
            10'b1011000011: o_power = 10'd 586;  // alpha^586
            10'b0110001111: o_power = 10'd 587;  // alpha^587
            10'b1100011110: o_power = 10'd 588;  // alpha^588
            10'b1000110101: o_power = 10'd 589;  // alpha^589
            10'b0001100011: o_power = 10'd 590;  // alpha^590
            10'b0011000110: o_power = 10'd 591;  // alpha^591
            10'b0110001100: o_power = 10'd 592;  // alpha^592
            10'b1100011000: o_power = 10'd 593;  // alpha^593
            10'b1000111001: o_power = 10'd 594;  // alpha^594
            10'b0001111011: o_power = 10'd 595;  // alpha^595
            10'b0011110110: o_power = 10'd 596;  // alpha^596
            10'b0111101100: o_power = 10'd 597;  // alpha^597
            10'b1111011000: o_power = 10'd 598;  // alpha^598
            10'b1110111001: o_power = 10'd 599;  // alpha^599
            10'b1101111011: o_power = 10'd 600;  // alpha^600
            10'b1011111111: o_power = 10'd 601;  // alpha^601
            10'b0111110111: o_power = 10'd 602;  // alpha^602
            10'b1111101110: o_power = 10'd 603;  // alpha^603
            10'b1111010101: o_power = 10'd 604;  // alpha^604
            10'b1110100011: o_power = 10'd 605;  // alpha^605
            10'b1101001111: o_power = 10'd 606;  // alpha^606
            10'b1010010111: o_power = 10'd 607;  // alpha^607
            10'b0100100111: o_power = 10'd 608;  // alpha^608
            10'b1001001110: o_power = 10'd 609;  // alpha^609
            10'b0010010101: o_power = 10'd 610;  // alpha^610
            10'b0100101010: o_power = 10'd 611;  // alpha^611
            10'b1001010100: o_power = 10'd 612;  // alpha^612
            10'b0010100001: o_power = 10'd 613;  // alpha^613
            10'b0101000010: o_power = 10'd 614;  // alpha^614
            10'b1010000100: o_power = 10'd 615;  // alpha^615
            10'b0100000001: o_power = 10'd 616;  // alpha^616
            10'b1000000010: o_power = 10'd 617;  // alpha^617
            10'b0000001101: o_power = 10'd 618;  // alpha^618
            10'b0000011010: o_power = 10'd 619;  // alpha^619
            10'b0000110100: o_power = 10'd 620;  // alpha^620
            10'b0001101000: o_power = 10'd 621;  // alpha^621
            10'b0011010000: o_power = 10'd 622;  // alpha^622
            10'b0110100000: o_power = 10'd 623;  // alpha^623
            10'b1101000000: o_power = 10'd 624;  // alpha^624
            10'b1010001001: o_power = 10'd 625;  // alpha^625
            10'b0100011011: o_power = 10'd 626;  // alpha^626
            10'b1000110110: o_power = 10'd 627;  // alpha^627
            10'b0001100101: o_power = 10'd 628;  // alpha^628
            10'b0011001010: o_power = 10'd 629;  // alpha^629
            10'b0110010100: o_power = 10'd 630;  // alpha^630
            10'b1100101000: o_power = 10'd 631;  // alpha^631
            10'b1001011001: o_power = 10'd 632;  // alpha^632
            10'b0010111011: o_power = 10'd 633;  // alpha^633
            10'b0101110110: o_power = 10'd 634;  // alpha^634
            10'b1011101100: o_power = 10'd 635;  // alpha^635
            10'b0111010001: o_power = 10'd 636;  // alpha^636
            10'b1110100010: o_power = 10'd 637;  // alpha^637
            10'b1101001101: o_power = 10'd 638;  // alpha^638
            10'b1010010011: o_power = 10'd 639;  // alpha^639
            10'b0100101111: o_power = 10'd 640;  // alpha^640
            10'b1001011110: o_power = 10'd 641;  // alpha^641
            10'b0010110101: o_power = 10'd 642;  // alpha^642
            10'b0101101010: o_power = 10'd 643;  // alpha^643
            10'b1011010100: o_power = 10'd 644;  // alpha^644
            10'b0110100001: o_power = 10'd 645;  // alpha^645
            10'b1101000010: o_power = 10'd 646;  // alpha^646
            10'b1010001101: o_power = 10'd 647;  // alpha^647
            10'b0100010011: o_power = 10'd 648;  // alpha^648
            10'b1000100110: o_power = 10'd 649;  // alpha^649
            10'b0001000101: o_power = 10'd 650;  // alpha^650
            10'b0010001010: o_power = 10'd 651;  // alpha^651
            10'b0100010100: o_power = 10'd 652;  // alpha^652
            10'b1000101000: o_power = 10'd 653;  // alpha^653
            10'b0001011001: o_power = 10'd 654;  // alpha^654
            10'b0010110010: o_power = 10'd 655;  // alpha^655
            10'b0101100100: o_power = 10'd 656;  // alpha^656
            10'b1011001000: o_power = 10'd 657;  // alpha^657
            10'b0110011001: o_power = 10'd 658;  // alpha^658
            10'b1100110010: o_power = 10'd 659;  // alpha^659
            10'b1001101101: o_power = 10'd 660;  // alpha^660
            10'b0011010011: o_power = 10'd 661;  // alpha^661
            10'b0110100110: o_power = 10'd 662;  // alpha^662
            10'b1101001100: o_power = 10'd 663;  // alpha^663
            10'b1010010001: o_power = 10'd 664;  // alpha^664
            10'b0100101011: o_power = 10'd 665;  // alpha^665
            10'b1001010110: o_power = 10'd 666;  // alpha^666
            10'b0010100101: o_power = 10'd 667;  // alpha^667
            10'b0101001010: o_power = 10'd 668;  // alpha^668
            10'b1010010100: o_power = 10'd 669;  // alpha^669
            10'b0100100001: o_power = 10'd 670;  // alpha^670
            10'b1001000010: o_power = 10'd 671;  // alpha^671
            10'b0010001101: o_power = 10'd 672;  // alpha^672
            10'b0100011010: o_power = 10'd 673;  // alpha^673
            10'b1000110100: o_power = 10'd 674;  // alpha^674
            10'b0001100001: o_power = 10'd 675;  // alpha^675
            10'b0011000010: o_power = 10'd 676;  // alpha^676
            10'b0110000100: o_power = 10'd 677;  // alpha^677
            10'b1100001000: o_power = 10'd 678;  // alpha^678
            10'b1000011001: o_power = 10'd 679;  // alpha^679
            10'b0000111011: o_power = 10'd 680;  // alpha^680
            10'b0001110110: o_power = 10'd 681;  // alpha^681
            10'b0011101100: o_power = 10'd 682;  // alpha^682
            10'b0111011000: o_power = 10'd 683;  // alpha^683
            10'b1110110000: o_power = 10'd 684;  // alpha^684
            10'b1101101001: o_power = 10'd 685;  // alpha^685
            10'b1011011011: o_power = 10'd 686;  // alpha^686
            10'b0110111111: o_power = 10'd 687;  // alpha^687
            10'b1101111110: o_power = 10'd 688;  // alpha^688
            10'b1011110101: o_power = 10'd 689;  // alpha^689
            10'b0111100011: o_power = 10'd 690;  // alpha^690
            10'b1111000110: o_power = 10'd 691;  // alpha^691
            10'b1110000101: o_power = 10'd 692;  // alpha^692
            10'b1100000011: o_power = 10'd 693;  // alpha^693
            10'b1000001111: o_power = 10'd 694;  // alpha^694
            10'b0000010111: o_power = 10'd 695;  // alpha^695
            10'b0000101110: o_power = 10'd 696;  // alpha^696
            10'b0001011100: o_power = 10'd 697;  // alpha^697
            10'b0010111000: o_power = 10'd 698;  // alpha^698
            10'b0101110000: o_power = 10'd 699;  // alpha^699
            10'b1011100000: o_power = 10'd 700;  // alpha^700
            10'b0111001001: o_power = 10'd 701;  // alpha^701
            10'b1110010010: o_power = 10'd 702;  // alpha^702
            10'b1100101101: o_power = 10'd 703;  // alpha^703
            10'b1001010011: o_power = 10'd 704;  // alpha^704
            10'b0010101111: o_power = 10'd 705;  // alpha^705
            10'b0101011110: o_power = 10'd 706;  // alpha^706
            10'b1010111100: o_power = 10'd 707;  // alpha^707
            10'b0101110001: o_power = 10'd 708;  // alpha^708
            10'b1011100010: o_power = 10'd 709;  // alpha^709
            10'b0111001101: o_power = 10'd 710;  // alpha^710
            10'b1110011010: o_power = 10'd 711;  // alpha^711
            10'b1100111101: o_power = 10'd 712;  // alpha^712
            10'b1001110011: o_power = 10'd 713;  // alpha^713
            10'b0011101111: o_power = 10'd 714;  // alpha^714
            10'b0111011110: o_power = 10'd 715;  // alpha^715
            10'b1110111100: o_power = 10'd 716;  // alpha^716
            10'b1101110001: o_power = 10'd 717;  // alpha^717
            10'b1011101011: o_power = 10'd 718;  // alpha^718
            10'b0111011111: o_power = 10'd 719;  // alpha^719
            10'b1110111110: o_power = 10'd 720;  // alpha^720
            10'b1101110101: o_power = 10'd 721;  // alpha^721
            10'b1011100011: o_power = 10'd 722;  // alpha^722
            10'b0111001111: o_power = 10'd 723;  // alpha^723
            10'b1110011110: o_power = 10'd 724;  // alpha^724
            10'b1100110101: o_power = 10'd 725;  // alpha^725
            10'b1001100011: o_power = 10'd 726;  // alpha^726
            10'b0011001111: o_power = 10'd 727;  // alpha^727
            10'b0110011110: o_power = 10'd 728;  // alpha^728
            10'b1100111100: o_power = 10'd 729;  // alpha^729
            10'b1001110001: o_power = 10'd 730;  // alpha^730
            10'b0011101011: o_power = 10'd 731;  // alpha^731
            10'b0111010110: o_power = 10'd 732;  // alpha^732
            10'b1110101100: o_power = 10'd 733;  // alpha^733
            10'b1101010001: o_power = 10'd 734;  // alpha^734
            10'b1010101011: o_power = 10'd 735;  // alpha^735
            10'b0101011111: o_power = 10'd 736;  // alpha^736
            10'b1010111110: o_power = 10'd 737;  // alpha^737
            10'b0101110101: o_power = 10'd 738;  // alpha^738
            10'b1011101010: o_power = 10'd 739;  // alpha^739
            10'b0111011101: o_power = 10'd 740;  // alpha^740
            10'b1110111010: o_power = 10'd 741;  // alpha^741
            10'b1101111101: o_power = 10'd 742;  // alpha^742
            10'b1011110011: o_power = 10'd 743;  // alpha^743
            10'b0111101111: o_power = 10'd 744;  // alpha^744
            10'b1111011110: o_power = 10'd 745;  // alpha^745
            10'b1110110101: o_power = 10'd 746;  // alpha^746
            10'b1101100011: o_power = 10'd 747;  // alpha^747
            10'b1011001111: o_power = 10'd 748;  // alpha^748
            10'b0110010111: o_power = 10'd 749;  // alpha^749
            10'b1100101110: o_power = 10'd 750;  // alpha^750
            10'b1001010101: o_power = 10'd 751;  // alpha^751
            10'b0010100011: o_power = 10'd 752;  // alpha^752
            10'b0101000110: o_power = 10'd 753;  // alpha^753
            10'b1010001100: o_power = 10'd 754;  // alpha^754
            10'b0100010001: o_power = 10'd 755;  // alpha^755
            10'b1000100010: o_power = 10'd 756;  // alpha^756
            10'b0001001101: o_power = 10'd 757;  // alpha^757
            10'b0010011010: o_power = 10'd 758;  // alpha^758
            10'b0100110100: o_power = 10'd 759;  // alpha^759
            10'b1001101000: o_power = 10'd 760;  // alpha^760
            10'b0011011001: o_power = 10'd 761;  // alpha^761
            10'b0110110010: o_power = 10'd 762;  // alpha^762
            10'b1101100100: o_power = 10'd 763;  // alpha^763
            10'b1011000001: o_power = 10'd 764;  // alpha^764
            10'b0110001011: o_power = 10'd 765;  // alpha^765
            10'b1100010110: o_power = 10'd 766;  // alpha^766
            10'b1000100101: o_power = 10'd 767;  // alpha^767
            10'b0001000011: o_power = 10'd 768;  // alpha^768
            10'b0010000110: o_power = 10'd 769;  // alpha^769
            10'b0100001100: o_power = 10'd 770;  // alpha^770
            10'b1000011000: o_power = 10'd 771;  // alpha^771
            10'b0000111001: o_power = 10'd 772;  // alpha^772
            10'b0001110010: o_power = 10'd 773;  // alpha^773
            10'b0011100100: o_power = 10'd 774;  // alpha^774
            10'b0111001000: o_power = 10'd 775;  // alpha^775
            10'b1110010000: o_power = 10'd 776;  // alpha^776
            10'b1100101001: o_power = 10'd 777;  // alpha^777
            10'b1001011011: o_power = 10'd 778;  // alpha^778
            10'b0010111111: o_power = 10'd 779;  // alpha^779
            10'b0101111110: o_power = 10'd 780;  // alpha^780
            10'b1011111100: o_power = 10'd 781;  // alpha^781
            10'b0111110001: o_power = 10'd 782;  // alpha^782
            10'b1111100010: o_power = 10'd 783;  // alpha^783
            10'b1111001101: o_power = 10'd 784;  // alpha^784
            10'b1110010011: o_power = 10'd 785;  // alpha^785
            10'b1100101111: o_power = 10'd 786;  // alpha^786
            10'b1001010111: o_power = 10'd 787;  // alpha^787
            10'b0010100111: o_power = 10'd 788;  // alpha^788
            10'b0101001110: o_power = 10'd 789;  // alpha^789
            10'b1010011100: o_power = 10'd 790;  // alpha^790
            10'b0100110001: o_power = 10'd 791;  // alpha^791
            10'b1001100010: o_power = 10'd 792;  // alpha^792
            10'b0011001101: o_power = 10'd 793;  // alpha^793
            10'b0110011010: o_power = 10'd 794;  // alpha^794
            10'b1100110100: o_power = 10'd 795;  // alpha^795
            10'b1001100001: o_power = 10'd 796;  // alpha^796
            10'b0011001011: o_power = 10'd 797;  // alpha^797
            10'b0110010110: o_power = 10'd 798;  // alpha^798
            10'b1100101100: o_power = 10'd 799;  // alpha^799
            10'b1001010001: o_power = 10'd 800;  // alpha^800
            10'b0010101011: o_power = 10'd 801;  // alpha^801
            10'b0101010110: o_power = 10'd 802;  // alpha^802
            10'b1010101100: o_power = 10'd 803;  // alpha^803
            10'b0101010001: o_power = 10'd 804;  // alpha^804
            10'b1010100010: o_power = 10'd 805;  // alpha^805
            10'b0101001101: o_power = 10'd 806;  // alpha^806
            10'b1010011010: o_power = 10'd 807;  // alpha^807
            10'b0100111101: o_power = 10'd 808;  // alpha^808
            10'b1001111010: o_power = 10'd 809;  // alpha^809
            10'b0011111101: o_power = 10'd 810;  // alpha^810
            10'b0111111010: o_power = 10'd 811;  // alpha^811
            10'b1111110100: o_power = 10'd 812;  // alpha^812
            10'b1111100001: o_power = 10'd 813;  // alpha^813
            10'b1111001011: o_power = 10'd 814;  // alpha^814
            10'b1110011111: o_power = 10'd 815;  // alpha^815
            10'b1100110111: o_power = 10'd 816;  // alpha^816
            10'b1001100111: o_power = 10'd 817;  // alpha^817
            10'b0011000111: o_power = 10'd 818;  // alpha^818
            10'b0110001110: o_power = 10'd 819;  // alpha^819
            10'b1100011100: o_power = 10'd 820;  // alpha^820
            10'b1000110001: o_power = 10'd 821;  // alpha^821
            10'b0001101011: o_power = 10'd 822;  // alpha^822
            10'b0011010110: o_power = 10'd 823;  // alpha^823
            10'b0110101100: o_power = 10'd 824;  // alpha^824
            10'b1101011000: o_power = 10'd 825;  // alpha^825
            10'b1010111001: o_power = 10'd 826;  // alpha^826
            10'b0101111011: o_power = 10'd 827;  // alpha^827
            10'b1011110110: o_power = 10'd 828;  // alpha^828
            10'b0111100101: o_power = 10'd 829;  // alpha^829
            10'b1111001010: o_power = 10'd 830;  // alpha^830
            10'b1110011101: o_power = 10'd 831;  // alpha^831
            10'b1100110011: o_power = 10'd 832;  // alpha^832
            10'b1001101111: o_power = 10'd 833;  // alpha^833
            10'b0011010111: o_power = 10'd 834;  // alpha^834
            10'b0110101110: o_power = 10'd 835;  // alpha^835
            10'b1101011100: o_power = 10'd 836;  // alpha^836
            10'b1010110001: o_power = 10'd 837;  // alpha^837
            10'b0101101011: o_power = 10'd 838;  // alpha^838
            10'b1011010110: o_power = 10'd 839;  // alpha^839
            10'b0110100101: o_power = 10'd 840;  // alpha^840
            10'b1101001010: o_power = 10'd 841;  // alpha^841
            10'b1010011101: o_power = 10'd 842;  // alpha^842
            10'b0100110011: o_power = 10'd 843;  // alpha^843
            10'b1001100110: o_power = 10'd 844;  // alpha^844
            10'b0011000101: o_power = 10'd 845;  // alpha^845
            10'b0110001010: o_power = 10'd 846;  // alpha^846
            10'b1100010100: o_power = 10'd 847;  // alpha^847
            10'b1000100001: o_power = 10'd 848;  // alpha^848
            10'b0001001011: o_power = 10'd 849;  // alpha^849
            10'b0010010110: o_power = 10'd 850;  // alpha^850
            10'b0100101100: o_power = 10'd 851;  // alpha^851
            10'b1001011000: o_power = 10'd 852;  // alpha^852
            10'b0010111001: o_power = 10'd 853;  // alpha^853
            10'b0101110010: o_power = 10'd 854;  // alpha^854
            10'b1011100100: o_power = 10'd 855;  // alpha^855
            10'b0111000001: o_power = 10'd 856;  // alpha^856
            10'b1110000010: o_power = 10'd 857;  // alpha^857
            10'b1100001101: o_power = 10'd 858;  // alpha^858
            10'b1000010011: o_power = 10'd 859;  // alpha^859
            10'b0000101111: o_power = 10'd 860;  // alpha^860
            10'b0001011110: o_power = 10'd 861;  // alpha^861
            10'b0010111100: o_power = 10'd 862;  // alpha^862
            10'b0101111000: o_power = 10'd 863;  // alpha^863
            10'b1011110000: o_power = 10'd 864;  // alpha^864
            10'b0111101001: o_power = 10'd 865;  // alpha^865
            10'b1111010010: o_power = 10'd 866;  // alpha^866
            10'b1110101101: o_power = 10'd 867;  // alpha^867
            10'b1101010011: o_power = 10'd 868;  // alpha^868
            10'b1010101111: o_power = 10'd 869;  // alpha^869
            10'b0101010111: o_power = 10'd 870;  // alpha^870
            10'b1010101110: o_power = 10'd 871;  // alpha^871
            10'b0101010101: o_power = 10'd 872;  // alpha^872
            10'b1010101010: o_power = 10'd 873;  // alpha^873
            10'b0101011101: o_power = 10'd 874;  // alpha^874
            10'b1010111010: o_power = 10'd 875;  // alpha^875
            10'b0101111101: o_power = 10'd 876;  // alpha^876
            10'b1011111010: o_power = 10'd 877;  // alpha^877
            10'b0111111101: o_power = 10'd 878;  // alpha^878
            10'b1111111010: o_power = 10'd 879;  // alpha^879
            10'b1111111101: o_power = 10'd 880;  // alpha^880
            10'b1111110011: o_power = 10'd 881;  // alpha^881
            10'b1111101111: o_power = 10'd 882;  // alpha^882
            10'b1111010111: o_power = 10'd 883;  // alpha^883
            10'b1110100111: o_power = 10'd 884;  // alpha^884
            10'b1101000111: o_power = 10'd 885;  // alpha^885
            10'b1010000111: o_power = 10'd 886;  // alpha^886
            10'b0100000111: o_power = 10'd 887;  // alpha^887
            10'b1000001110: o_power = 10'd 888;  // alpha^888
            10'b0000010101: o_power = 10'd 889;  // alpha^889
            10'b0000101010: o_power = 10'd 890;  // alpha^890
            10'b0001010100: o_power = 10'd 891;  // alpha^891
            10'b0010101000: o_power = 10'd 892;  // alpha^892
            10'b0101010000: o_power = 10'd 893;  // alpha^893
            10'b1010100000: o_power = 10'd 894;  // alpha^894
            10'b0101001001: o_power = 10'd 895;  // alpha^895
            10'b1010010010: o_power = 10'd 896;  // alpha^896
            10'b0100101101: o_power = 10'd 897;  // alpha^897
            10'b1001011010: o_power = 10'd 898;  // alpha^898
            10'b0010111101: o_power = 10'd 899;  // alpha^899
            10'b0101111010: o_power = 10'd 900;  // alpha^900
            10'b1011110100: o_power = 10'd 901;  // alpha^901
            10'b0111100001: o_power = 10'd 902;  // alpha^902
            10'b1111000010: o_power = 10'd 903;  // alpha^903
            10'b1110001101: o_power = 10'd 904;  // alpha^904
            10'b1100010011: o_power = 10'd 905;  // alpha^905
            10'b1000101111: o_power = 10'd 906;  // alpha^906
            10'b0001010111: o_power = 10'd 907;  // alpha^907
            10'b0010101110: o_power = 10'd 908;  // alpha^908
            10'b0101011100: o_power = 10'd 909;  // alpha^909
            10'b1010111000: o_power = 10'd 910;  // alpha^910
            10'b0101111001: o_power = 10'd 911;  // alpha^911
            10'b1011110010: o_power = 10'd 912;  // alpha^912
            10'b0111101101: o_power = 10'd 913;  // alpha^913
            10'b1111011010: o_power = 10'd 914;  // alpha^914
            10'b1110111101: o_power = 10'd 915;  // alpha^915
            10'b1101110011: o_power = 10'd 916;  // alpha^916
            10'b1011101111: o_power = 10'd 917;  // alpha^917
            10'b0111010111: o_power = 10'd 918;  // alpha^918
            10'b1110101110: o_power = 10'd 919;  // alpha^919
            10'b1101010101: o_power = 10'd 920;  // alpha^920
            10'b1010100011: o_power = 10'd 921;  // alpha^921
            10'b0101001111: o_power = 10'd 922;  // alpha^922
            10'b1010011110: o_power = 10'd 923;  // alpha^923
            10'b0100110101: o_power = 10'd 924;  // alpha^924
            10'b1001101010: o_power = 10'd 925;  // alpha^925
            10'b0011011101: o_power = 10'd 926;  // alpha^926
            10'b0110111010: o_power = 10'd 927;  // alpha^927
            10'b1101110100: o_power = 10'd 928;  // alpha^928
            10'b1011100001: o_power = 10'd 929;  // alpha^929
            10'b0111001011: o_power = 10'd 930;  // alpha^930
            10'b1110010110: o_power = 10'd 931;  // alpha^931
            10'b1100100101: o_power = 10'd 932;  // alpha^932
            10'b1001000011: o_power = 10'd 933;  // alpha^933
            10'b0010001111: o_power = 10'd 934;  // alpha^934
            10'b0100011110: o_power = 10'd 935;  // alpha^935
            10'b1000111100: o_power = 10'd 936;  // alpha^936
            10'b0001110001: o_power = 10'd 937;  // alpha^937
            10'b0011100010: o_power = 10'd 938;  // alpha^938
            10'b0111000100: o_power = 10'd 939;  // alpha^939
            10'b1110001000: o_power = 10'd 940;  // alpha^940
            10'b1100011001: o_power = 10'd 941;  // alpha^941
            10'b1000111011: o_power = 10'd 942;  // alpha^942
            10'b0001111111: o_power = 10'd 943;  // alpha^943
            10'b0011111110: o_power = 10'd 944;  // alpha^944
            10'b0111111100: o_power = 10'd 945;  // alpha^945
            10'b1111111000: o_power = 10'd 946;  // alpha^946
            10'b1111111001: o_power = 10'd 947;  // alpha^947
            10'b1111111011: o_power = 10'd 948;  // alpha^948
            10'b1111111111: o_power = 10'd 949;  // alpha^949
            10'b1111110111: o_power = 10'd 950;  // alpha^950
            10'b1111100111: o_power = 10'd 951;  // alpha^951
            10'b1111000111: o_power = 10'd 952;  // alpha^952
            10'b1110000111: o_power = 10'd 953;  // alpha^953
            10'b1100000111: o_power = 10'd 954;  // alpha^954
            10'b1000000111: o_power = 10'd 955;  // alpha^955
            10'b0000000111: o_power = 10'd 956;  // alpha^956
            10'b0000001110: o_power = 10'd 957;  // alpha^957
            10'b0000011100: o_power = 10'd 958;  // alpha^958
            10'b0000111000: o_power = 10'd 959;  // alpha^959
            10'b0001110000: o_power = 10'd 960;  // alpha^960
            10'b0011100000: o_power = 10'd 961;  // alpha^961
            10'b0111000000: o_power = 10'd 962;  // alpha^962
            10'b1110000000: o_power = 10'd 963;  // alpha^963
            10'b1100001001: o_power = 10'd 964;  // alpha^964
            10'b1000011011: o_power = 10'd 965;  // alpha^965
            10'b0000111111: o_power = 10'd 966;  // alpha^966
            10'b0001111110: o_power = 10'd 967;  // alpha^967
            10'b0011111100: o_power = 10'd 968;  // alpha^968
            10'b0111111000: o_power = 10'd 969;  // alpha^969
            10'b1111110000: o_power = 10'd 970;  // alpha^970
            10'b1111101001: o_power = 10'd 971;  // alpha^971
            10'b1111011011: o_power = 10'd 972;  // alpha^972
            10'b1110111111: o_power = 10'd 973;  // alpha^973
            10'b1101110111: o_power = 10'd 974;  // alpha^974
            10'b1011100111: o_power = 10'd 975;  // alpha^975
            10'b0111000111: o_power = 10'd 976;  // alpha^976
            10'b1110001110: o_power = 10'd 977;  // alpha^977
            10'b1100010101: o_power = 10'd 978;  // alpha^978
            10'b1000100011: o_power = 10'd 979;  // alpha^979
            10'b0001001111: o_power = 10'd 980;  // alpha^980
            10'b0010011110: o_power = 10'd 981;  // alpha^981
            10'b0100111100: o_power = 10'd 982;  // alpha^982
            10'b1001111000: o_power = 10'd 983;  // alpha^983
            10'b0011111001: o_power = 10'd 984;  // alpha^984
            10'b0111110010: o_power = 10'd 985;  // alpha^985
            10'b1111100100: o_power = 10'd 986;  // alpha^986
            10'b1111000001: o_power = 10'd 987;  // alpha^987
            10'b1110001011: o_power = 10'd 988;  // alpha^988
            10'b1100011111: o_power = 10'd 989;  // alpha^989
            10'b1000110111: o_power = 10'd 990;  // alpha^990
            10'b0001100111: o_power = 10'd 991;  // alpha^991
            10'b0011001110: o_power = 10'd 992;  // alpha^992
            10'b0110011100: o_power = 10'd 993;  // alpha^993
            10'b1100111000: o_power = 10'd 994;  // alpha^994
            10'b1001111001: o_power = 10'd 995;  // alpha^995
            10'b0011111011: o_power = 10'd 996;  // alpha^996
            10'b0111110110: o_power = 10'd 997;  // alpha^997
            10'b1111101100: o_power = 10'd 998;  // alpha^998
            10'b1111010001: o_power = 10'd 999;  // alpha^999
            10'b1110101011: o_power = 10'd1000;  // alpha^1000
            10'b1101011111: o_power = 10'd1001;  // alpha^1001
            10'b1010110111: o_power = 10'd1002;  // alpha^1002
            10'b0101100111: o_power = 10'd1003;  // alpha^1003
            10'b1011001110: o_power = 10'd1004;  // alpha^1004
            10'b0110010101: o_power = 10'd1005;  // alpha^1005
            10'b1100101010: o_power = 10'd1006;  // alpha^1006
            10'b1001011101: o_power = 10'd1007;  // alpha^1007
            10'b0010110011: o_power = 10'd1008;  // alpha^1008
            10'b0101100110: o_power = 10'd1009;  // alpha^1009
            10'b1011001100: o_power = 10'd1010;  // alpha^1010
            10'b0110010001: o_power = 10'd1011;  // alpha^1011
            10'b1100100010: o_power = 10'd1012;  // alpha^1012
            10'b1001001101: o_power = 10'd1013;  // alpha^1013
            10'b0010010011: o_power = 10'd1014;  // alpha^1014
            10'b0100100110: o_power = 10'd1015;  // alpha^1015
            10'b1001001100: o_power = 10'd1016;  // alpha^1016
            10'b0010010001: o_power = 10'd1017;  // alpha^1017
            10'b0100100010: o_power = 10'd1018;  // alpha^1018
            10'b1001000100: o_power = 10'd1019;  // alpha^1019
            10'b0010000001: o_power = 10'd1020;  // alpha^1020
            10'b0100000010: o_power = 10'd1021;  // alpha^1021
            10'b1000000100: o_power = 10'd1022;  // alpha^1022
        endcase
    end

endmodule