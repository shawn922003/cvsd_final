module chien_search(
    
);

endmodule