module flip_alpha(
    input i_clk,
    input i_rst_n,

    input [63:0] i_data,

    input i_code,

    input i_clear,
    input i_wen,

    output [9:0] o_alpha1,
    output [9:0] o_alpha2,

    output [9:0] o_p1,
    output [9:0] o_p2,

    output o_valid
);


endmodule